----------------------------------------------------------
--  sim_cfg.vhd
--		Configuration for ZX97 simulation
--		=================================
--
--  04/24/97	Bodo Wenzel	Creation
--  11/14/97	Bodo Wenzel	Some polish
----------------------------------------------------------

-- the configuration (very simple!) ----------------------

configuration simu of tb is
  for beh
  end for;
end;

-- end ---------------------------------------------------
