library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ROM81hll is
	port(
		Clk	: in std_logic;
		AIn	: in std_logic_vector(11 downto 0);
		D	: out std_logic_vector(7 downto 0)
	);
end ROM81hll;

architecture rtl of ROM81hll is
	signal A	: std_logic_vector(12 downto 0);
begin
	A(12 downto 10) <= "100";
	process (Clk)
	begin
		if Clk'event and Clk = '1' then
			A(9 downto 0) <= AIn(9 downto 0);
		end if;
	end process;
	process (A)
	begin
		case to_integer(unsigned(A)) is
		when 004096 => D <= "10011010";	-- 0x1000
		when 004097 => D <= "00001101";	-- 0x1001
		when 004098 => D <= "11010110";	-- 0x1002
		when 004099 => D <= "11000100";	-- 0x1003
		when 004100 => D <= "00111000";	-- 0x1004
		when 004101 => D <= "11111001";	-- 0x1005
		when 004102 => D <= "00000001";	-- 0x1006
		when 004103 => D <= "11101100";	-- 0x1007
		when 004104 => D <= "00000100";	-- 0x1008
		when 004105 => D <= "11111110";	-- 0x1009
		when 004106 => D <= "00010011";	-- 0x100A
		when 004107 => D <= "00101000";	-- 0x100B
		when 004108 => D <= "00010011";	-- 0x100C
		when 004109 => D <= "00110000";	-- 0x100D
		when 004110 => D <= "11110000";	-- 0x100E
		when 004111 => D <= "00000110";	-- 0x100F
		when 004112 => D <= "00010000";	-- 0x1010
		when 004113 => D <= "11000110";	-- 0x1011
		when 004114 => D <= "11011001";	-- 0x1012
		when 004115 => D <= "01001111";	-- 0x1013
		when 004116 => D <= "11111110";	-- 0x1014
		when 004117 => D <= "11011100";	-- 0x1015
		when 004118 => D <= "00110000";	-- 0x1016
		when 004119 => D <= "00000010";	-- 0x1017
		when 004120 => D <= "11001011";	-- 0x1018
		when 004121 => D <= "10110001";	-- 0x1019
		when 004122 => D <= "11111110";	-- 0x101A
		when 004123 => D <= "11101010";	-- 0x101B
		when 004124 => D <= "00111000";	-- 0x101C
		when 004125 => D <= "00000010";	-- 0x101D
		when 004126 => D <= "11001011";	-- 0x101E
		when 004127 => D <= "10111001";	-- 0x101F
		when 004128 => D <= "11000101";	-- 0x1020
		when 004129 => D <= "11100111";	-- 0x1021
		when 004130 => D <= "11000011";	-- 0x1022
		when 004131 => D <= "01011001";	-- 0x1023
		when 004132 => D <= "00001111";	-- 0x1024
		when 004133 => D <= "11111110";	-- 0x1025
		when 004134 => D <= "00100110";	-- 0x1026
		when 004135 => D <= "00111000";	-- 0x1027
		when 004136 => D <= "00011110";	-- 0x1028
		when 004137 => D <= "11001101";	-- 0x1029
		when 004138 => D <= "00011100";	-- 0x102A
		when 004139 => D <= "00010001";	-- 0x102B
		when 004140 => D <= "11011010";	-- 0x102C
		when 004141 => D <= "01001011";	-- 0x102D
		when 004142 => D <= "00001101";	-- 0x102E
		when 004143 => D <= "11001100";	-- 0x102F
		when 004144 => D <= "10100111";	-- 0x1030
		when 004145 => D <= "00010001";	-- 0x1031
		when 004146 => D <= "00111010";	-- 0x1032
		when 004147 => D <= "00000001";	-- 0x1033
		when 004148 => D <= "01000000";	-- 0x1034
		when 004149 => D <= "11111110";	-- 0x1035
		when 004150 => D <= "11000000";	-- 0x1036
		when 004151 => D <= "00111000";	-- 0x1037
		when 004152 => D <= "01001110";	-- 0x1038
		when 004153 => D <= "00100011";	-- 0x1039
		when 004154 => D <= "11101101";	-- 0x103A
		when 004155 => D <= "01011011";	-- 0x103B
		when 004156 => D <= "00011100";	-- 0x103C
		when 004157 => D <= "01000000";	-- 0x103D
		when 004158 => D <= "11001101";	-- 0x103E
		when 004159 => D <= "11110110";	-- 0x103F
		when 004160 => D <= "00011001";	-- 0x1040
		when 004161 => D <= "11101011";	-- 0x1041
		when 004162 => D <= "00100010";	-- 0x1042
		when 004163 => D <= "00011100";	-- 0x1043
		when 004164 => D <= "01000000";	-- 0x1044
		when 004165 => D <= "00011000";	-- 0x1045
		when 004166 => D <= "01000000";	-- 0x1046
		when 004167 => D <= "11001101";	-- 0x1047
		when 004168 => D <= "10100110";	-- 0x1048
		when 004169 => D <= "00001101";	-- 0x1049
		when 004170 => D <= "00100000";	-- 0x104A
		when 004171 => D <= "00100011";	-- 0x104B
		when 004172 => D <= "11001101";	-- 0x104C
		when 004173 => D <= "11011001";	-- 0x104D
		when 004174 => D <= "00010100";	-- 0x104E
		when 004175 => D <= "11011111";	-- 0x104F
		when 004176 => D <= "00000001";	-- 0x1050
		when 004177 => D <= "00000110";	-- 0x1051
		when 004178 => D <= "00000000";	-- 0x1052
		when 004179 => D <= "11001101";	-- 0x1053
		when 004180 => D <= "10011110";	-- 0x1054
		when 004181 => D <= "00001001";	-- 0x1055
		when 004182 => D <= "00100011";	-- 0x1056
		when 004183 => D <= "00110110";	-- 0x1057
		when 004184 => D <= "01111110";	-- 0x1058
		when 004185 => D <= "00100011";	-- 0x1059
		when 004186 => D <= "11101011";	-- 0x105A
		when 004187 => D <= "00101010";	-- 0x105B
		when 004188 => D <= "00011100";	-- 0x105C
		when 004189 => D <= "01000000";	-- 0x105D
		when 004190 => D <= "00001110";	-- 0x105E
		when 004191 => D <= "00000101";	-- 0x105F
		when 004192 => D <= "10100111";	-- 0x1060
		when 004193 => D <= "11101101";	-- 0x1061
		when 004194 => D <= "01000010";	-- 0x1062
		when 004195 => D <= "00100010";	-- 0x1063
		when 004196 => D <= "00011100";	-- 0x1064
		when 004197 => D <= "01000000";	-- 0x1065
		when 004198 => D <= "11101101";	-- 0x1066
		when 004199 => D <= "10110000";	-- 0x1067
		when 004200 => D <= "11101011";	-- 0x1068
		when 004201 => D <= "00101011";	-- 0x1069
		when 004202 => D <= "11001101";	-- 0x106A
		when 004203 => D <= "01001100";	-- 0x106B
		when 004204 => D <= "00000000";	-- 0x106C
		when 004205 => D <= "00011000";	-- 0x106D
		when 004206 => D <= "00010100";	-- 0x106E
		when 004207 => D <= "11100111";	-- 0x106F
		when 004208 => D <= "11111110";	-- 0x1070
		when 004209 => D <= "01111110";	-- 0x1071
		when 004210 => D <= "00100000";	-- 0x1072
		when 004211 => D <= "11111011";	-- 0x1073
		when 004212 => D <= "00100011";	-- 0x1074
		when 004213 => D <= "11101101";	-- 0x1075
		when 004214 => D <= "01011011";	-- 0x1076
		when 004215 => D <= "00011100";	-- 0x1077
		when 004216 => D <= "01000000";	-- 0x1078
		when 004217 => D <= "11001101";	-- 0x1079
		when 004218 => D <= "11110110";	-- 0x107A
		when 004219 => D <= "00011001";	-- 0x107B
		when 004220 => D <= "11101101";	-- 0x107C
		when 004221 => D <= "01010011";	-- 0x107D
		when 004222 => D <= "00011100";	-- 0x107E
		when 004223 => D <= "01000000";	-- 0x107F
		when 004224 => D <= "00100010";	-- 0x1080
		when 004225 => D <= "00010110";	-- 0x1081
		when 004226 => D <= "01000000";	-- 0x1082
		when 004227 => D <= "11111101";	-- 0x1083
		when 004228 => D <= "11001011";	-- 0x1084
		when 004229 => D <= "00000001";	-- 0x1085
		when 004230 => D <= "11110110";	-- 0x1086
		when 004231 => D <= "11011111";	-- 0x1087
		when 004232 => D <= "11111110";	-- 0x1088
		when 004233 => D <= "00010000";	-- 0x1089
		when 004234 => D <= "00100000";	-- 0x108A
		when 004235 => D <= "00001100";	-- 0x108B
		when 004236 => D <= "11111101";	-- 0x108C
		when 004237 => D <= "11001011";	-- 0x108D
		when 004238 => D <= "00000001";	-- 0x108E
		when 004239 => D <= "01110110";	-- 0x108F
		when 004240 => D <= "00100000";	-- 0x1090
		when 004241 => D <= "00101010";	-- 0x1091
		when 004242 => D <= "11001101";	-- 0x1092
		when 004243 => D <= "01100011";	-- 0x1093
		when 004244 => D <= "00010010";	-- 0x1094
		when 004245 => D <= "11100111";	-- 0x1095
		when 004246 => D <= "00011000";	-- 0x1096
		when 004247 => D <= "11110000";	-- 0x1097
		when 004248 => D <= "00000001";	-- 0x1098
		when 004249 => D <= "11000011";	-- 0x1099
		when 004250 => D <= "00000000";	-- 0x109A
		when 004251 => D <= "11111110";	-- 0x109B
		when 004252 => D <= "00010010";	-- 0x109C
		when 004253 => D <= "00111000";	-- 0x109D
		when 004254 => D <= "00011101";	-- 0x109E
		when 004255 => D <= "11010110";	-- 0x109F
		when 004256 => D <= "00010110";	-- 0x10A0
		when 004257 => D <= "00110000";	-- 0x10A1
		when 004258 => D <= "00000100";	-- 0x10A2
		when 004259 => D <= "11000110";	-- 0x10A3
		when 004260 => D <= "00001101";	-- 0x10A4
		when 004261 => D <= "00011000";	-- 0x10A5
		when 004262 => D <= "00001110";	-- 0x10A6
		when 004263 => D <= "11111110";	-- 0x10A7
		when 004264 => D <= "00000011";	-- 0x10A8
		when 004265 => D <= "00111000";	-- 0x10A9
		when 004266 => D <= "00001010";	-- 0x10AA
		when 004267 => D <= "11010110";	-- 0x10AB
		when 004268 => D <= "11000010";	-- 0x10AC
		when 004269 => D <= "00111000";	-- 0x10AD
		when 004270 => D <= "00001101";	-- 0x10AE
		when 004271 => D <= "11111110";	-- 0x10AF
		when 004272 => D <= "00000110";	-- 0x10B0
		when 004273 => D <= "00110000";	-- 0x10B1
		when 004274 => D <= "00001001";	-- 0x10B2
		when 004275 => D <= "11000110";	-- 0x10B3
		when 004276 => D <= "00000011";	-- 0x10B4
		when 004277 => D <= "10000001";	-- 0x10B5
		when 004278 => D <= "01001111";	-- 0x10B6
		when 004279 => D <= "00100001";	-- 0x10B7
		when 004280 => D <= "01001100";	-- 0x10B8
		when 004281 => D <= "00010000";	-- 0x10B9
		when 004282 => D <= "00001001";	-- 0x10BA
		when 004283 => D <= "01000110";	-- 0x10BB
		when 004284 => D <= "11010001";	-- 0x10BC
		when 004285 => D <= "01111010";	-- 0x10BD
		when 004286 => D <= "10111000";	-- 0x10BE
		when 004287 => D <= "00111000";	-- 0x10BF
		when 004288 => D <= "00101100";	-- 0x10C0
		when 004289 => D <= "10100111";	-- 0x10C1
		when 004290 => D <= "11001010";	-- 0x10C2
		when 004291 => D <= "00011000";	-- 0x10C3
		when 004292 => D <= "00000000";	-- 0x10C4
		when 004293 => D <= "11000101";	-- 0x10C5
		when 004294 => D <= "11010101";	-- 0x10C6
		when 004295 => D <= "11001101";	-- 0x10C7
		when 004296 => D <= "10100110";	-- 0x10C8
		when 004297 => D <= "00001101";	-- 0x10C9
		when 004298 => D <= "00101000";	-- 0x10CA
		when 004299 => D <= "00001001";	-- 0x10CB
		when 004300 => D <= "01111011";	-- 0x10CC
		when 004301 => D <= "11100110";	-- 0x10CD
		when 004302 => D <= "00111111";	-- 0x10CE
		when 004303 => D <= "01000111";	-- 0x10CF
		when 004304 => D <= "11101111";	-- 0x10D0
		when 004305 => D <= "00110111";	-- 0x10D1
		when 004306 => D <= "00110100";	-- 0x10D2
		when 004307 => D <= "00011000";	-- 0x10D3
		when 004308 => D <= "00001001";	-- 0x10D4
		when 004309 => D <= "01111011";	-- 0x10D5
		when 004310 => D <= "11111101";	-- 0x10D6
		when 004311 => D <= "10101110";	-- 0x10D7
		when 004312 => D <= "00000001";	-- 0x10D8
		when 004313 => D <= "11100110";	-- 0x10D9
		when 004314 => D <= "01000000";	-- 0x10DA
		when 004315 => D <= "11000010";	-- 0x10DB
		when 004316 => D <= "10011010";	-- 0x10DC
		when 004317 => D <= "00001101";	-- 0x10DD
		when 004318 => D <= "11010001";	-- 0x10DE
		when 004319 => D <= "00100001";	-- 0x10DF
		when 004320 => D <= "00000001";	-- 0x10E0
		when 004321 => D <= "01000000";	-- 0x10E1
		when 004322 => D <= "11001011";	-- 0x10E2
		when 004323 => D <= "11110110";	-- 0x10E3
		when 004324 => D <= "11001011";	-- 0x10E4
		when 004325 => D <= "01111011";	-- 0x10E5
		when 004326 => D <= "00100000";	-- 0x10E6
		when 004327 => D <= "00000010";	-- 0x10E7
		when 004328 => D <= "11001011";	-- 0x10E8
		when 004329 => D <= "10110110";	-- 0x10E9
		when 004330 => D <= "11000001";	-- 0x10EA
		when 004331 => D <= "00011000";	-- 0x10EB
		when 004332 => D <= "11001111";	-- 0x10EC
		when 004333 => D <= "11010101";	-- 0x10ED
		when 004334 => D <= "01111001";	-- 0x10EE
		when 004335 => D <= "11111101";	-- 0x10EF
		when 004336 => D <= "11001011";	-- 0x10F0
		when 004337 => D <= "00000001";	-- 0x10F1
		when 004338 => D <= "01110110";	-- 0x10F2
		when 004339 => D <= "00100000";	-- 0x10F3
		when 004340 => D <= "00010101";	-- 0x10F4
		when 004341 => D <= "11100110";	-- 0x10F5
		when 004342 => D <= "00111111";	-- 0x10F6
		when 004343 => D <= "11000110";	-- 0x10F7
		when 004344 => D <= "00001000";	-- 0x10F8
		when 004345 => D <= "01001111";	-- 0x10F9
		when 004346 => D <= "11111110";	-- 0x10FA
		when 004347 => D <= "00010000";	-- 0x10FB
		when 004348 => D <= "00100000";	-- 0x10FC
		when 004349 => D <= "00000100";	-- 0x10FD
		when 004350 => D <= "11001011";	-- 0x10FE
		when 004351 => D <= "11110001";	-- 0x10FF
		when 004352 => D <= "00011000";	-- 0x1100
		when 004353 => D <= "00001000";	-- 0x1101
		when 004354 => D <= "00111000";	-- 0x1102
		when 004355 => D <= "11010111";	-- 0x1103
		when 004356 => D <= "11111110";	-- 0x1104
		when 004357 => D <= "00010111";	-- 0x1105
		when 004358 => D <= "00101000";	-- 0x1106
		when 004359 => D <= "00000010";	-- 0x1107
		when 004360 => D <= "11001011";	-- 0x1108
		when 004361 => D <= "11111001";	-- 0x1109
		when 004362 => D <= "11000101";	-- 0x110A
		when 004363 => D <= "11100111";	-- 0x110B
		when 004364 => D <= "11000011";	-- 0x110C
		when 004365 => D <= "01011001";	-- 0x110D
		when 004366 => D <= "00001111";	-- 0x110E
		when 004367 => D <= "00000110";	-- 0x110F
		when 004368 => D <= "00001000";	-- 0x1110
		when 004369 => D <= "00001000";	-- 0x1111
		when 004370 => D <= "00001010";	-- 0x1112
		when 004371 => D <= "00000010";	-- 0x1113
		when 004372 => D <= "00000011";	-- 0x1114
		when 004373 => D <= "00000101";	-- 0x1115
		when 004374 => D <= "00000101";	-- 0x1116
		when 004375 => D <= "00000101";	-- 0x1117
		when 004376 => D <= "00000101";	-- 0x1118
		when 004377 => D <= "00000101";	-- 0x1119
		when 004378 => D <= "00000101";	-- 0x111A
		when 004379 => D <= "00000110";	-- 0x111B
		when 004380 => D <= "11111101";	-- 0x111C
		when 004381 => D <= "11001011";	-- 0x111D
		when 004382 => D <= "00000001";	-- 0x111E
		when 004383 => D <= "11110110";	-- 0x111F
		when 004384 => D <= "11011111";	-- 0x1120
		when 004385 => D <= "11001101";	-- 0x1121
		when 004386 => D <= "11001110";	-- 0x1122
		when 004387 => D <= "00010100";	-- 0x1123
		when 004388 => D <= "11010010";	-- 0x1124
		when 004389 => D <= "10011010";	-- 0x1125
		when 004390 => D <= "00001101";	-- 0x1126
		when 004391 => D <= "11100101";	-- 0x1127
		when 004392 => D <= "01001111";	-- 0x1128
		when 004393 => D <= "11100111";	-- 0x1129
		when 004394 => D <= "11100101";	-- 0x112A
		when 004395 => D <= "11001011";	-- 0x112B
		when 004396 => D <= "10101001";	-- 0x112C
		when 004397 => D <= "11111110";	-- 0x112D
		when 004398 => D <= "00010000";	-- 0x112E
		when 004399 => D <= "00101000";	-- 0x112F
		when 004400 => D <= "00010111";	-- 0x1130
		when 004401 => D <= "11001011";	-- 0x1131
		when 004402 => D <= "11110001";	-- 0x1132
		when 004403 => D <= "11111110";	-- 0x1133
		when 004404 => D <= "00001101";	-- 0x1134
		when 004405 => D <= "00101000";	-- 0x1135
		when 004406 => D <= "00001100";	-- 0x1136
		when 004407 => D <= "11001011";	-- 0x1137
		when 004408 => D <= "11101001";	-- 0x1138
		when 004409 => D <= "11001101";	-- 0x1139
		when 004410 => D <= "11010010";	-- 0x113A
		when 004411 => D <= "00010100";	-- 0x113B
		when 004412 => D <= "00110000";	-- 0x113C
		when 004413 => D <= "00001010";	-- 0x113D
		when 004414 => D <= "11001011";	-- 0x113E
		when 004415 => D <= "10110001";	-- 0x113F
		when 004416 => D <= "11100111";	-- 0x1140
		when 004417 => D <= "00011000";	-- 0x1141
		when 004418 => D <= "11110110";	-- 0x1142
		when 004419 => D <= "11100111";	-- 0x1143
		when 004420 => D <= "11111101";	-- 0x1144
		when 004421 => D <= "11001011";	-- 0x1145
		when 004422 => D <= "00000001";	-- 0x1146
		when 004423 => D <= "10110110";	-- 0x1147
		when 004424 => D <= "01000001";	-- 0x1148
		when 004425 => D <= "11001101";	-- 0x1149
		when 004426 => D <= "10100110";	-- 0x114A
		when 004427 => D <= "00001101";	-- 0x114B
		when 004428 => D <= "00100000";	-- 0x114C
		when 004429 => D <= "00001000";	-- 0x114D
		when 004430 => D <= "01111001";	-- 0x114E
		when 004431 => D <= "11100110";	-- 0x114F
		when 004432 => D <= "11100000";	-- 0x1150
		when 004433 => D <= "11001011";	-- 0x1151
		when 004434 => D <= "11111111";	-- 0x1152
		when 004435 => D <= "01001111";	-- 0x1153
		when 004436 => D <= "00011000";	-- 0x1154
		when 004437 => D <= "00110100";	-- 0x1155
		when 004438 => D <= "00101010";	-- 0x1156
		when 004439 => D <= "00010000";	-- 0x1157
		when 004440 => D <= "01000000";	-- 0x1158
		when 004441 => D <= "01111110";	-- 0x1159
		when 004442 => D <= "11100110";	-- 0x115A
		when 004443 => D <= "01111111";	-- 0x115B
		when 004444 => D <= "00101000";	-- 0x115C
		when 004445 => D <= "00101010";	-- 0x115D
		when 004446 => D <= "10111001";	-- 0x115E
		when 004447 => D <= "00100000";	-- 0x115F
		when 004448 => D <= "00011111";	-- 0x1160
		when 004449 => D <= "00010111";	-- 0x1161
		when 004450 => D <= "10000111";	-- 0x1162
		when 004451 => D <= "11110010";	-- 0x1163
		when 004452 => D <= "10010101";	-- 0x1164
		when 004453 => D <= "00010001";	-- 0x1165
		when 004454 => D <= "00111000";	-- 0x1166
		when 004455 => D <= "00101101";	-- 0x1167
		when 004456 => D <= "11010001";	-- 0x1168
		when 004457 => D <= "11010101";	-- 0x1169
		when 004458 => D <= "11100101";	-- 0x116A
		when 004459 => D <= "00100011";	-- 0x116B
		when 004460 => D <= "00011010";	-- 0x116C
		when 004461 => D <= "00010011";	-- 0x116D
		when 004462 => D <= "10100111";	-- 0x116E
		when 004463 => D <= "00101000";	-- 0x116F
		when 004464 => D <= "11111011";	-- 0x1170
		when 004465 => D <= "10111110";	-- 0x1171
		when 004466 => D <= "00101000";	-- 0x1172
		when 004467 => D <= "11110111";	-- 0x1173
		when 004468 => D <= "11110110";	-- 0x1174
		when 004469 => D <= "10000000";	-- 0x1175
		when 004470 => D <= "10111110";	-- 0x1176
		when 004471 => D <= "00100000";	-- 0x1177
		when 004472 => D <= "00000110";	-- 0x1178
		when 004473 => D <= "00011010";	-- 0x1179
		when 004474 => D <= "11001101";	-- 0x117A
		when 004475 => D <= "11010010";	-- 0x117B
		when 004476 => D <= "00010100";	-- 0x117C
		when 004477 => D <= "00110000";	-- 0x117D
		when 004478 => D <= "00010101";	-- 0x117E
		when 004479 => D <= "11100001";	-- 0x117F
		when 004480 => D <= "11000101";	-- 0x1180
		when 004481 => D <= "11001101";	-- 0x1181
		when 004482 => D <= "11110010";	-- 0x1182
		when 004483 => D <= "00001001";	-- 0x1183
		when 004484 => D <= "11101011";	-- 0x1184
		when 004485 => D <= "11000001";	-- 0x1185
		when 004486 => D <= "00011000";	-- 0x1186
		when 004487 => D <= "11010001";	-- 0x1187
		when 004488 => D <= "11001011";	-- 0x1188
		when 004489 => D <= "11111000";	-- 0x1189
		when 004490 => D <= "11010001";	-- 0x118A
		when 004491 => D <= "11011111";	-- 0x118B
		when 004492 => D <= "11111110";	-- 0x118C
		when 004493 => D <= "00010000";	-- 0x118D
		when 004494 => D <= "00101000";	-- 0x118E
		when 004495 => D <= "00001001";	-- 0x118F
		when 004496 => D <= "11001011";	-- 0x1190
		when 004497 => D <= "11101000";	-- 0x1191
		when 004498 => D <= "00011000";	-- 0x1192
		when 004499 => D <= "00001101";	-- 0x1193
		when 004500 => D <= "11010001";	-- 0x1194
		when 004501 => D <= "11010001";	-- 0x1195
		when 004502 => D <= "11010001";	-- 0x1196
		when 004503 => D <= "11100101";	-- 0x1197
		when 004504 => D <= "11011111";	-- 0x1198
		when 004505 => D <= "11001101";	-- 0x1199
		when 004506 => D <= "11010010";	-- 0x119A
		when 004507 => D <= "00010100";	-- 0x119B
		when 004508 => D <= "00110000";	-- 0x119C
		when 004509 => D <= "00000011";	-- 0x119D
		when 004510 => D <= "11100111";	-- 0x119E
		when 004511 => D <= "00011000";	-- 0x119F
		when 004512 => D <= "11111000";	-- 0x11A0
		when 004513 => D <= "11100001";	-- 0x11A1
		when 004514 => D <= "11001011";	-- 0x11A2
		when 004515 => D <= "00010000";	-- 0x11A3
		when 004516 => D <= "11001011";	-- 0x11A4
		when 004517 => D <= "01110000";	-- 0x11A5
		when 004518 => D <= "11001001";	-- 0x11A6
		when 004519 => D <= "10101111";	-- 0x11A7
		when 004520 => D <= "01000111";	-- 0x11A8
		when 004521 => D <= "11001011";	-- 0x11A9
		when 004522 => D <= "01111001";	-- 0x11AA
		when 004523 => D <= "00100000";	-- 0x11AB
		when 004524 => D <= "01001011";	-- 0x11AC
		when 004525 => D <= "11001011";	-- 0x11AD
		when 004526 => D <= "01111110";	-- 0x11AE
		when 004527 => D <= "00100000";	-- 0x11AF
		when 004528 => D <= "00001110";	-- 0x11B0
		when 004529 => D <= "00111100";	-- 0x11B1
		when 004530 => D <= "00100011";	-- 0x11B2
		when 004531 => D <= "01001110";	-- 0x11B3
		when 004532 => D <= "00100011";	-- 0x11B4
		when 004533 => D <= "01000110";	-- 0x11B5
		when 004534 => D <= "00100011";	-- 0x11B6
		when 004535 => D <= "11101011";	-- 0x11B7
		when 004536 => D <= "11001101";	-- 0x11B8
		when 004537 => D <= "11000011";	-- 0x11B9
		when 004538 => D <= "00010010";	-- 0x11BA
		when 004539 => D <= "11011111";	-- 0x11BB
		when 004540 => D <= "11000011";	-- 0x11BC
		when 004541 => D <= "01011010";	-- 0x11BD
		when 004542 => D <= "00010010";	-- 0x11BE
		when 004543 => D <= "00100011";	-- 0x11BF
		when 004544 => D <= "00100011";	-- 0x11C0
		when 004545 => D <= "00100011";	-- 0x11C1
		when 004546 => D <= "01000110";	-- 0x11C2
		when 004547 => D <= "11001011";	-- 0x11C3
		when 004548 => D <= "01110001";	-- 0x11C4
		when 004549 => D <= "00101000";	-- 0x11C5
		when 004550 => D <= "00001010";	-- 0x11C6
		when 004551 => D <= "00000101";	-- 0x11C7
		when 004552 => D <= "00101000";	-- 0x11C8
		when 004553 => D <= "11101000";	-- 0x11C9
		when 004554 => D <= "11101011";	-- 0x11CA
		when 004555 => D <= "11011111";	-- 0x11CB
		when 004556 => D <= "11111110";	-- 0x11CC
		when 004557 => D <= "00010000";	-- 0x11CD
		when 004558 => D <= "00100000";	-- 0x11CE
		when 004559 => D <= "01100001";	-- 0x11CF
		when 004560 => D <= "11101011";	-- 0x11D0
		when 004561 => D <= "11101011";	-- 0x11D1
		when 004562 => D <= "00011000";	-- 0x11D2
		when 004563 => D <= "00100100";	-- 0x11D3
		when 004564 => D <= "11100101";	-- 0x11D4
		when 004565 => D <= "11011111";	-- 0x11D5
		when 004566 => D <= "11100001";	-- 0x11D6
		when 004567 => D <= "11111110";	-- 0x11D7
		when 004568 => D <= "00011010";	-- 0x11D8
		when 004569 => D <= "00101000";	-- 0x11D9
		when 004570 => D <= "00100000";	-- 0x11DA
		when 004571 => D <= "11001011";	-- 0x11DB
		when 004572 => D <= "01111001";	-- 0x11DC
		when 004573 => D <= "00101000";	-- 0x11DD
		when 004574 => D <= "01010010";	-- 0x11DE
		when 004575 => D <= "11001011";	-- 0x11DF
		when 004576 => D <= "01110001";	-- 0x11E0
		when 004577 => D <= "00100000";	-- 0x11E1
		when 004578 => D <= "00000110";	-- 0x11E2
		when 004579 => D <= "11111110";	-- 0x11E3
		when 004580 => D <= "00010001";	-- 0x11E4
		when 004581 => D <= "00100000";	-- 0x11E5
		when 004582 => D <= "00111100";	-- 0x11E6
		when 004583 => D <= "11100111";	-- 0x11E7
		when 004584 => D <= "11001001";	-- 0x11E8
		when 004585 => D <= "11111110";	-- 0x11E9
		when 004586 => D <= "00010001";	-- 0x11EA
		when 004587 => D <= "00101000";	-- 0x11EB
		when 004588 => D <= "01101100";	-- 0x11EC
		when 004589 => D <= "11111110";	-- 0x11ED
		when 004590 => D <= "11011111";	-- 0x11EE
		when 004591 => D <= "00100000";	-- 0x11EF
		when 004592 => D <= "00110010";	-- 0x11F0
		when 004593 => D <= "11011111";	-- 0x11F1
		when 004594 => D <= "00101011";	-- 0x11F2
		when 004595 => D <= "00100010";	-- 0x11F3
		when 004596 => D <= "00010110";	-- 0x11F4
		when 004597 => D <= "01000000";	-- 0x11F5
		when 004598 => D <= "00011000";	-- 0x11F6
		when 004599 => D <= "01011110";	-- 0x11F7
		when 004600 => D <= "00100001";	-- 0x11F8
		when 004601 => D <= "00000000";	-- 0x11F9
		when 004602 => D <= "00000000";	-- 0x11FA
		when 004603 => D <= "11100101";	-- 0x11FB
		when 004604 => D <= "11100111";	-- 0x11FC
		when 004605 => D <= "11100001";	-- 0x11FD
		when 004606 => D <= "01111001";	-- 0x11FE
		when 004607 => D <= "11111110";	-- 0x11FF
		when 004608 => D <= "11000000";	-- 0x1200
		when 004609 => D <= "00100000";	-- 0x1201
		when 004610 => D <= "00001001";	-- 0x1202
		when 004611 => D <= "11011111";	-- 0x1203
		when 004612 => D <= "11111110";	-- 0x1204
		when 004613 => D <= "00010001";	-- 0x1205
		when 004614 => D <= "00101000";	-- 0x1206
		when 004615 => D <= "01010001";	-- 0x1207
		when 004616 => D <= "11111110";	-- 0x1208
		when 004617 => D <= "11011111";	-- 0x1209
		when 004618 => D <= "00101000";	-- 0x120A
		when 004619 => D <= "11100101";	-- 0x120B
		when 004620 => D <= "11000101";	-- 0x120C
		when 004621 => D <= "11100101";	-- 0x120D
		when 004622 => D <= "11001101";	-- 0x120E
		when 004623 => D <= "11111111";	-- 0x120F
		when 004624 => D <= "00010010";	-- 0x1210
		when 004625 => D <= "11100011";	-- 0x1211
		when 004626 => D <= "11101011";	-- 0x1212
		when 004627 => D <= "11001101";	-- 0x1213
		when 004628 => D <= "11011101";	-- 0x1214
		when 004629 => D <= "00010010";	-- 0x1215
		when 004630 => D <= "00111000";	-- 0x1216
		when 004631 => D <= "00011001";	-- 0x1217
		when 004632 => D <= "00001011";	-- 0x1218
		when 004633 => D <= "11001101";	-- 0x1219
		when 004634 => D <= "00000101";	-- 0x121A
		when 004635 => D <= "00010011";	-- 0x121B
		when 004636 => D <= "00001001";	-- 0x121C
		when 004637 => D <= "11010001";	-- 0x121D
		when 004638 => D <= "11000001";	-- 0x121E
		when 004639 => D <= "00010000";	-- 0x121F
		when 004640 => D <= "10110011";	-- 0x1220
		when 004641 => D <= "11001011";	-- 0x1221
		when 004642 => D <= "01111001";	-- 0x1222
		when 004643 => D <= "00100000";	-- 0x1223
		when 004644 => D <= "01100110";	-- 0x1224
		when 004645 => D <= "11100101";	-- 0x1225
		when 004646 => D <= "11001011";	-- 0x1226
		when 004647 => D <= "01110001";	-- 0x1227
		when 004648 => D <= "00100000";	-- 0x1228
		when 004649 => D <= "00010011";	-- 0x1229
		when 004650 => D <= "01000010";	-- 0x122A
		when 004651 => D <= "01001011";	-- 0x122B
		when 004652 => D <= "11011111";	-- 0x122C
		when 004653 => D <= "11111110";	-- 0x122D
		when 004654 => D <= "00010001";	-- 0x122E
		when 004655 => D <= "00101000";	-- 0x122F
		when 004656 => D <= "00000010";	-- 0x1230
		when 004657 => D <= "11001111";	-- 0x1231
		when 004658 => D <= "00000010";	-- 0x1232
		when 004659 => D <= "11100111";	-- 0x1233
		when 004660 => D <= "11100001";	-- 0x1234
		when 004661 => D <= "00010001";	-- 0x1235
		when 004662 => D <= "00000101";	-- 0x1236
		when 004663 => D <= "00000000";	-- 0x1237
		when 004664 => D <= "11001101";	-- 0x1238
		when 004665 => D <= "00000101";	-- 0x1239
		when 004666 => D <= "00010011";	-- 0x123A
		when 004667 => D <= "00001001";	-- 0x123B
		when 004668 => D <= "11001001";	-- 0x123C
		when 004669 => D <= "11001101";	-- 0x123D
		when 004670 => D <= "11111111";	-- 0x123E
		when 004671 => D <= "00010010";	-- 0x123F
		when 004672 => D <= "11100011";	-- 0x1240
		when 004673 => D <= "11001101";	-- 0x1241
		when 004674 => D <= "00000101";	-- 0x1242
		when 004675 => D <= "00010011";	-- 0x1243
		when 004676 => D <= "11000001";	-- 0x1244
		when 004677 => D <= "00001001";	-- 0x1245
		when 004678 => D <= "00100011";	-- 0x1246
		when 004679 => D <= "01000010";	-- 0x1247
		when 004680 => D <= "01001011";	-- 0x1248
		when 004681 => D <= "11101011";	-- 0x1249
		when 004682 => D <= "11001101";	-- 0x124A
		when 004683 => D <= "11000010";	-- 0x124B
		when 004684 => D <= "00010010";	-- 0x124C
		when 004685 => D <= "11011111";	-- 0x124D
		when 004686 => D <= "11111110";	-- 0x124E
		when 004687 => D <= "00010001";	-- 0x124F
		when 004688 => D <= "00101000";	-- 0x1250
		when 004689 => D <= "00000111";	-- 0x1251
		when 004690 => D <= "11111110";	-- 0x1252
		when 004691 => D <= "00011010";	-- 0x1253
		when 004692 => D <= "00100000";	-- 0x1254
		when 004693 => D <= "11011011";	-- 0x1255
		when 004694 => D <= "11001101";	-- 0x1256
		when 004695 => D <= "01100011";	-- 0x1257
		when 004696 => D <= "00010010";	-- 0x1258
		when 004697 => D <= "11100111";	-- 0x1259
		when 004698 => D <= "11111110";	-- 0x125A
		when 004699 => D <= "00010000";	-- 0x125B
		when 004700 => D <= "00101000";	-- 0x125C
		when 004701 => D <= "11111000";	-- 0x125D
		when 004702 => D <= "11111101";	-- 0x125E
		when 004703 => D <= "11001011";	-- 0x125F
		when 004704 => D <= "00000001";	-- 0x1260
		when 004705 => D <= "10110110";	-- 0x1261
		when 004706 => D <= "11001001";	-- 0x1262
		when 004707 => D <= "11001101";	-- 0x1263
		when 004708 => D <= "10100110";	-- 0x1264
		when 004709 => D <= "00001101";	-- 0x1265
		when 004710 => D <= "11000100";	-- 0x1266
		when 004711 => D <= "11111000";	-- 0x1267
		when 004712 => D <= "00010011";	-- 0x1268
		when 004713 => D <= "11100111";	-- 0x1269
		when 004714 => D <= "11111110";	-- 0x126A
		when 004715 => D <= "00010001";	-- 0x126B
		when 004716 => D <= "00101000";	-- 0x126C
		when 004717 => D <= "01010000";	-- 0x126D
		when 004718 => D <= "11010101";	-- 0x126E
		when 004719 => D <= "10101111";	-- 0x126F
		when 004720 => D <= "11110101";	-- 0x1270
		when 004721 => D <= "11000101";	-- 0x1271
		when 004722 => D <= "00010001";	-- 0x1272
		when 004723 => D <= "00000001";	-- 0x1273
		when 004724 => D <= "00000000";	-- 0x1274
		when 004725 => D <= "11011111";	-- 0x1275
		when 004726 => D <= "11100001";	-- 0x1276
		when 004727 => D <= "11111110";	-- 0x1277
		when 004728 => D <= "11011111";	-- 0x1278
		when 004729 => D <= "00101000";	-- 0x1279
		when 004730 => D <= "00010111";	-- 0x127A
		when 004731 => D <= "11110001";	-- 0x127B
		when 004732 => D <= "11001101";	-- 0x127C
		when 004733 => D <= "11011110";	-- 0x127D
		when 004734 => D <= "00010010";	-- 0x127E
		when 004735 => D <= "11110101";	-- 0x127F
		when 004736 => D <= "01010000";	-- 0x1280
		when 004737 => D <= "01011001";	-- 0x1281
		when 004738 => D <= "11100101";	-- 0x1282
		when 004739 => D <= "11011111";	-- 0x1283
		when 004740 => D <= "11100001";	-- 0x1284
		when 004741 => D <= "11111110";	-- 0x1285
		when 004742 => D <= "11011111";	-- 0x1286
		when 004743 => D <= "00101000";	-- 0x1287
		when 004744 => D <= "00001001";	-- 0x1288
		when 004745 => D <= "11111110";	-- 0x1289
		when 004746 => D <= "00010001";	-- 0x128A
		when 004747 => D <= "11000010";	-- 0x128B
		when 004748 => D <= "10011010";	-- 0x128C
		when 004749 => D <= "00001101";	-- 0x128D
		when 004750 => D <= "01100010";	-- 0x128E
		when 004751 => D <= "01101011";	-- 0x128F
		when 004752 => D <= "00011000";	-- 0x1290
		when 004753 => D <= "00010011";	-- 0x1291
		when 004754 => D <= "11100101";	-- 0x1292
		when 004755 => D <= "11100111";	-- 0x1293
		when 004756 => D <= "11100001";	-- 0x1294
		when 004757 => D <= "11111110";	-- 0x1295
		when 004758 => D <= "00010001";	-- 0x1296
		when 004759 => D <= "00101000";	-- 0x1297
		when 004760 => D <= "00001100";	-- 0x1298
		when 004761 => D <= "11110001";	-- 0x1299
		when 004762 => D <= "11001101";	-- 0x129A
		when 004763 => D <= "11011110";	-- 0x129B
		when 004764 => D <= "00010010";	-- 0x129C
		when 004765 => D <= "11110101";	-- 0x129D
		when 004766 => D <= "11011111";	-- 0x129E
		when 004767 => D <= "01100000";	-- 0x129F
		when 004768 => D <= "01101001";	-- 0x12A0
		when 004769 => D <= "11111110";	-- 0x12A1
		when 004770 => D <= "00010001";	-- 0x12A2
		when 004771 => D <= "00100000";	-- 0x12A3
		when 004772 => D <= "11100110";	-- 0x12A4
		when 004773 => D <= "11110001";	-- 0x12A5
		when 004774 => D <= "11100011";	-- 0x12A6
		when 004775 => D <= "00011001";	-- 0x12A7
		when 004776 => D <= "00101011";	-- 0x12A8
		when 004777 => D <= "11100011";	-- 0x12A9
		when 004778 => D <= "10100111";	-- 0x12AA
		when 004779 => D <= "11101101";	-- 0x12AB
		when 004780 => D <= "01010010";	-- 0x12AC
		when 004781 => D <= "00000001";	-- 0x12AD
		when 004782 => D <= "00000000";	-- 0x12AE
		when 004783 => D <= "00000000";	-- 0x12AF
		when 004784 => D <= "00111000";	-- 0x12B0
		when 004785 => D <= "00000111";	-- 0x12B1
		when 004786 => D <= "00100011";	-- 0x12B2
		when 004787 => D <= "10100111";	-- 0x12B3
		when 004788 => D <= "11111010";	-- 0x12B4
		when 004789 => D <= "00110001";	-- 0x12B5
		when 004790 => D <= "00010010";	-- 0x12B6
		when 004791 => D <= "01000100";	-- 0x12B7
		when 004792 => D <= "01001101";	-- 0x12B8
		when 004793 => D <= "11010001";	-- 0x12B9
		when 004794 => D <= "11111101";	-- 0x12BA
		when 004795 => D <= "11001011";	-- 0x12BB
		when 004796 => D <= "00000001";	-- 0x12BC
		when 004797 => D <= "10110110";	-- 0x12BD
		when 004798 => D <= "11001101";	-- 0x12BE
		when 004799 => D <= "10100110";	-- 0x12BF
		when 004800 => D <= "00001101";	-- 0x12C0
		when 004801 => D <= "11001000";	-- 0x12C1
		when 004802 => D <= "10101111";	-- 0x12C2
		when 004803 => D <= "11000101";	-- 0x12C3
		when 004804 => D <= "11001101";	-- 0x12C4
		when 004805 => D <= "11101011";	-- 0x12C5
		when 004806 => D <= "00011001";	-- 0x12C6
		when 004807 => D <= "11000001";	-- 0x12C7
		when 004808 => D <= "00101010";	-- 0x12C8
		when 004809 => D <= "00011100";	-- 0x12C9
		when 004810 => D <= "01000000";	-- 0x12CA
		when 004811 => D <= "01110111";	-- 0x12CB
		when 004812 => D <= "00100011";	-- 0x12CC
		when 004813 => D <= "01110011";	-- 0x12CD
		when 004814 => D <= "00100011";	-- 0x12CE
		when 004815 => D <= "01110010";	-- 0x12CF
		when 004816 => D <= "00100011";	-- 0x12D0
		when 004817 => D <= "01110001";	-- 0x12D1
		when 004818 => D <= "00100011";	-- 0x12D2
		when 004819 => D <= "01110000";	-- 0x12D3
		when 004820 => D <= "00100011";	-- 0x12D4
		when 004821 => D <= "00100010";	-- 0x12D5
		when 004822 => D <= "00011100";	-- 0x12D6
		when 004823 => D <= "01000000";	-- 0x12D7
		when 004824 => D <= "11111101";	-- 0x12D8
		when 004825 => D <= "11001011";	-- 0x12D9
		when 004826 => D <= "00000001";	-- 0x12DA
		when 004827 => D <= "10110110";	-- 0x12DB
		when 004828 => D <= "11001001";	-- 0x12DC
		when 004829 => D <= "10101111";	-- 0x12DD
		when 004830 => D <= "11010101";	-- 0x12DE
		when 004831 => D <= "11100101";	-- 0x12DF
		when 004832 => D <= "11110101";	-- 0x12E0
		when 004833 => D <= "11001101";	-- 0x12E1
		when 004834 => D <= "10010010";	-- 0x12E2
		when 004835 => D <= "00001101";	-- 0x12E3
		when 004836 => D <= "11110001";	-- 0x12E4
		when 004837 => D <= "11001101";	-- 0x12E5
		when 004838 => D <= "10100110";	-- 0x12E6
		when 004839 => D <= "00001101";	-- 0x12E7
		when 004840 => D <= "00101000";	-- 0x12E8
		when 004841 => D <= "00010010";	-- 0x12E9
		when 004842 => D <= "11110101";	-- 0x12EA
		when 004843 => D <= "11001101";	-- 0x12EB
		when 004844 => D <= "10100111";	-- 0x12EC
		when 004845 => D <= "00001110";	-- 0x12ED
		when 004846 => D <= "11010001";	-- 0x12EE
		when 004847 => D <= "01111000";	-- 0x12EF
		when 004848 => D <= "10110001";	-- 0x12F0
		when 004849 => D <= "00110111";	-- 0x12F1
		when 004850 => D <= "00101000";	-- 0x12F2
		when 004851 => D <= "00000101";	-- 0x12F3
		when 004852 => D <= "11100001";	-- 0x12F4
		when 004853 => D <= "11100101";	-- 0x12F5
		when 004854 => D <= "10100111";	-- 0x12F6
		when 004855 => D <= "11101101";	-- 0x12F7
		when 004856 => D <= "01000010";	-- 0x12F8
		when 004857 => D <= "01111010";	-- 0x12F9
		when 004858 => D <= "11011110";	-- 0x12FA
		when 004859 => D <= "00000000";	-- 0x12FB
		when 004860 => D <= "11100001";	-- 0x12FC
		when 004861 => D <= "11010001";	-- 0x12FD
		when 004862 => D <= "11001001";	-- 0x12FE
		when 004863 => D <= "11101011";	-- 0x12FF
		when 004864 => D <= "00100011";	-- 0x1300
		when 004865 => D <= "01011110";	-- 0x1301
		when 004866 => D <= "00100011";	-- 0x1302
		when 004867 => D <= "01010110";	-- 0x1303
		when 004868 => D <= "11001001";	-- 0x1304
		when 004869 => D <= "11001101";	-- 0x1305
		when 004870 => D <= "10100110";	-- 0x1306
		when 004871 => D <= "00001101";	-- 0x1307
		when 004872 => D <= "11001000";	-- 0x1308
		when 004873 => D <= "11000101";	-- 0x1309
		when 004874 => D <= "00000110";	-- 0x130A
		when 004875 => D <= "00010000";	-- 0x130B
		when 004876 => D <= "01111100";	-- 0x130C
		when 004877 => D <= "01001101";	-- 0x130D
		when 004878 => D <= "00100001";	-- 0x130E
		when 004879 => D <= "00000000";	-- 0x130F
		when 004880 => D <= "00000000";	-- 0x1310
		when 004881 => D <= "00101001";	-- 0x1311
		when 004882 => D <= "00111000";	-- 0x1312
		when 004883 => D <= "00000110";	-- 0x1313
		when 004884 => D <= "11001011";	-- 0x1314
		when 004885 => D <= "00010001";	-- 0x1315
		when 004886 => D <= "00010111";	-- 0x1316
		when 004887 => D <= "00110000";	-- 0x1317
		when 004888 => D <= "00000100";	-- 0x1318
		when 004889 => D <= "00011001";	-- 0x1319
		when 004890 => D <= "11011010";	-- 0x131A
		when 004891 => D <= "11010011";	-- 0x131B
		when 004892 => D <= "00001110";	-- 0x131C
		when 004893 => D <= "00010000";	-- 0x131D
		when 004894 => D <= "11110010";	-- 0x131E
		when 004895 => D <= "11000001";	-- 0x131F
		when 004896 => D <= "11001001";	-- 0x1320
		when 004897 => D <= "00101010";	-- 0x1321
		when 004898 => D <= "00010010";	-- 0x1322
		when 004899 => D <= "01000000";	-- 0x1323
		when 004900 => D <= "11111101";	-- 0x1324
		when 004901 => D <= "11001011";	-- 0x1325
		when 004902 => D <= "00101101";	-- 0x1326
		when 004903 => D <= "01001110";	-- 0x1327
		when 004904 => D <= "00101000";	-- 0x1328
		when 004905 => D <= "01000100";	-- 0x1329
		when 004906 => D <= "00000001";	-- 0x132A
		when 004907 => D <= "00000101";	-- 0x132B
		when 004908 => D <= "00000000";	-- 0x132C
		when 004909 => D <= "00000011";	-- 0x132D
		when 004910 => D <= "00100011";	-- 0x132E
		when 004911 => D <= "01111110";	-- 0x132F
		when 004912 => D <= "10100111";	-- 0x1330
		when 004913 => D <= "00101000";	-- 0x1331
		when 004914 => D <= "11111011";	-- 0x1332
		when 004915 => D <= "11001101";	-- 0x1333
		when 004916 => D <= "11010010";	-- 0x1334
		when 004917 => D <= "00010100";	-- 0x1335
		when 004918 => D <= "00111000";	-- 0x1336
		when 004919 => D <= "11110101";	-- 0x1337
		when 004920 => D <= "11111110";	-- 0x1338
		when 004921 => D <= "00001101";	-- 0x1339
		when 004922 => D <= "11001010";	-- 0x133A
		when 004923 => D <= "11001000";	-- 0x133B
		when 004924 => D <= "00010011";	-- 0x133C
		when 004925 => D <= "11110111";	-- 0x133D
		when 004926 => D <= "11010101";	-- 0x133E
		when 004927 => D <= "00101010";	-- 0x133F
		when 004928 => D <= "00010010";	-- 0x1340
		when 004929 => D <= "01000000";	-- 0x1341
		when 004930 => D <= "00011011";	-- 0x1342
		when 004931 => D <= "01111001";	-- 0x1343
		when 004932 => D <= "11010110";	-- 0x1344
		when 004933 => D <= "00000110";	-- 0x1345
		when 004934 => D <= "01000111";	-- 0x1346
		when 004935 => D <= "00111110";	-- 0x1347
		when 004936 => D <= "01000000";	-- 0x1348
		when 004937 => D <= "00101000";	-- 0x1349
		when 004938 => D <= "00001110";	-- 0x134A
		when 004939 => D <= "00100011";	-- 0x134B
		when 004940 => D <= "01111110";	-- 0x134C
		when 004941 => D <= "10100111";	-- 0x134D
		when 004942 => D <= "00101000";	-- 0x134E
		when 004943 => D <= "11111011";	-- 0x134F
		when 004944 => D <= "00010011";	-- 0x1350
		when 004945 => D <= "00010010";	-- 0x1351
		when 004946 => D <= "00010000";	-- 0x1352
		when 004947 => D <= "11110111";	-- 0x1353
		when 004948 => D <= "11110110";	-- 0x1354
		when 004949 => D <= "10000000";	-- 0x1355
		when 004950 => D <= "00010010";	-- 0x1356
		when 004951 => D <= "00111110";	-- 0x1357
		when 004952 => D <= "10000000";	-- 0x1358
		when 004953 => D <= "00101010";	-- 0x1359
		when 004954 => D <= "00010010";	-- 0x135A
		when 004955 => D <= "01000000";	-- 0x135B
		when 004956 => D <= "10101110";	-- 0x135C
		when 004957 => D <= "11100001";	-- 0x135D
		when 004958 => D <= "11001101";	-- 0x135E
		when 004959 => D <= "11100111";	-- 0x135F
		when 004960 => D <= "00010011";	-- 0x1360
		when 004961 => D <= "11100101";	-- 0x1361
		when 004962 => D <= "11101111";	-- 0x1362
		when 004963 => D <= "00000010";	-- 0x1363
		when 004964 => D <= "00110100";	-- 0x1364
		when 004965 => D <= "11100001";	-- 0x1365
		when 004966 => D <= "00000001";	-- 0x1366
		when 004967 => D <= "00000101";	-- 0x1367
		when 004968 => D <= "00000000";	-- 0x1368
		when 004969 => D <= "10100111";	-- 0x1369
		when 004970 => D <= "11101101";	-- 0x136A
		when 004971 => D <= "01000010";	-- 0x136B
		when 004972 => D <= "00011000";	-- 0x136C
		when 004973 => D <= "01000000";	-- 0x136D
		when 004974 => D <= "11111101";	-- 0x136E
		when 004975 => D <= "11001011";	-- 0x136F
		when 004976 => D <= "00000001";	-- 0x1370
		when 004977 => D <= "01110110";	-- 0x1371
		when 004978 => D <= "00101000";	-- 0x1372
		when 004979 => D <= "00000110";	-- 0x1373
		when 004980 => D <= "00010001";	-- 0x1374
		when 004981 => D <= "00000110";	-- 0x1375
		when 004982 => D <= "00000000";	-- 0x1376
		when 004983 => D <= "00011001";	-- 0x1377
		when 004984 => D <= "00011000";	-- 0x1378
		when 004985 => D <= "11100111";	-- 0x1379
		when 004986 => D <= "00101010";	-- 0x137A
		when 004987 => D <= "00010010";	-- 0x137B
		when 004988 => D <= "01000000";	-- 0x137C
		when 004989 => D <= "11101101";	-- 0x137D
		when 004990 => D <= "01001011";	-- 0x137E
		when 004991 => D <= "00101110";	-- 0x137F
		when 004992 => D <= "01000000";	-- 0x1380
		when 004993 => D <= "11111101";	-- 0x1381
		when 004994 => D <= "11001011";	-- 0x1382
		when 004995 => D <= "00101101";	-- 0x1383
		when 004996 => D <= "01000110";	-- 0x1384
		when 004997 => D <= "00100000";	-- 0x1385
		when 004998 => D <= "00110000";	-- 0x1386
		when 004999 => D <= "01111000";	-- 0x1387
		when 005000 => D <= "10110001";	-- 0x1388
		when 005001 => D <= "11001000";	-- 0x1389
		when 005002 => D <= "11100101";	-- 0x138A
		when 005003 => D <= "11110111";	-- 0x138B
		when 005004 => D <= "11010101";	-- 0x138C
		when 005005 => D <= "11000101";	-- 0x138D
		when 005006 => D <= "01010100";	-- 0x138E
		when 005007 => D <= "01011101";	-- 0x138F
		when 005008 => D <= "00100011";	-- 0x1390
		when 005009 => D <= "00110110";	-- 0x1391
		when 005010 => D <= "00000000";	-- 0x1392
		when 005011 => D <= "11101101";	-- 0x1393
		when 005012 => D <= "10111000";	-- 0x1394
		when 005013 => D <= "11100101";	-- 0x1395
		when 005014 => D <= "11001101";	-- 0x1396
		when 005015 => D <= "11111000";	-- 0x1397
		when 005016 => D <= "00010011";	-- 0x1398
		when 005017 => D <= "11100001";	-- 0x1399
		when 005018 => D <= "11100011";	-- 0x139A
		when 005019 => D <= "10100111";	-- 0x139B
		when 005020 => D <= "11101101";	-- 0x139C
		when 005021 => D <= "01000010";	-- 0x139D
		when 005022 => D <= "00001001";	-- 0x139E
		when 005023 => D <= "00110000";	-- 0x139F
		when 005024 => D <= "00000010";	-- 0x13A0
		when 005025 => D <= "01000100";	-- 0x13A1
		when 005026 => D <= "01001101";	-- 0x13A2
		when 005027 => D <= "11100011";	-- 0x13A3
		when 005028 => D <= "11101011";	-- 0x13A4
		when 005029 => D <= "01111000";	-- 0x13A5
		when 005030 => D <= "10110001";	-- 0x13A6
		when 005031 => D <= "00101000";	-- 0x13A7
		when 005032 => D <= "00000010";	-- 0x13A8
		when 005033 => D <= "11101101";	-- 0x13A9
		when 005034 => D <= "10110000";	-- 0x13AA
		when 005035 => D <= "11000001";	-- 0x13AB
		when 005036 => D <= "11010001";	-- 0x13AC
		when 005037 => D <= "11100001";	-- 0x13AD
		when 005038 => D <= "11101011";	-- 0x13AE
		when 005039 => D <= "01111000";	-- 0x13AF
		when 005040 => D <= "10110001";	-- 0x13B0
		when 005041 => D <= "11001000";	-- 0x13B1
		when 005042 => D <= "11010101";	-- 0x13B2
		when 005043 => D <= "11101101";	-- 0x13B3
		when 005044 => D <= "10110000";	-- 0x13B4
		when 005045 => D <= "11100001";	-- 0x13B5
		when 005046 => D <= "11001001";	-- 0x13B6
		when 005047 => D <= "00101011";	-- 0x13B7
		when 005048 => D <= "00101011";	-- 0x13B8
		when 005049 => D <= "00101011";	-- 0x13B9
		when 005050 => D <= "01111110";	-- 0x13BA
		when 005051 => D <= "11100101";	-- 0x13BB
		when 005052 => D <= "11000101";	-- 0x13BC
		when 005053 => D <= "11001101";	-- 0x13BD
		when 005054 => D <= "11001110";	-- 0x13BE
		when 005055 => D <= "00010011";	-- 0x13BF
		when 005056 => D <= "11000001";	-- 0x13C0
		when 005057 => D <= "11100001";	-- 0x13C1
		when 005058 => D <= "00000011";	-- 0x13C2
		when 005059 => D <= "00000011";	-- 0x13C3
		when 005060 => D <= "00000011";	-- 0x13C4
		when 005061 => D <= "11000011";	-- 0x13C5
		when 005062 => D <= "01100000";	-- 0x13C6
		when 005063 => D <= "00001010";	-- 0x13C7
		when 005064 => D <= "00111110";	-- 0x13C8
		when 005065 => D <= "01100000";	-- 0x13C9
		when 005066 => D <= "00101010";	-- 0x13CA
		when 005067 => D <= "00010010";	-- 0x13CB
		when 005068 => D <= "01000000";	-- 0x13CC
		when 005069 => D <= "10101110";	-- 0x13CD
		when 005070 => D <= "11110101";	-- 0x13CE
		when 005071 => D <= "11001101";	-- 0x13CF
		when 005072 => D <= "11111000";	-- 0x13D0
		when 005073 => D <= "00010011";	-- 0x13D1
		when 005074 => D <= "11101011";	-- 0x13D2
		when 005075 => D <= "00001001";	-- 0x13D3
		when 005076 => D <= "11100101";	-- 0x13D4
		when 005077 => D <= "00000011";	-- 0x13D5
		when 005078 => D <= "00000011";	-- 0x13D6
		when 005079 => D <= "00000011";	-- 0x13D7
		when 005080 => D <= "11110111";	-- 0x13D8
		when 005081 => D <= "11101011";	-- 0x13D9
		when 005082 => D <= "11100001";	-- 0x13DA
		when 005083 => D <= "00001011";	-- 0x13DB
		when 005084 => D <= "00001011";	-- 0x13DC
		when 005085 => D <= "11000101";	-- 0x13DD
		when 005086 => D <= "11101101";	-- 0x13DE
		when 005087 => D <= "10111000";	-- 0x13DF
		when 005088 => D <= "11101011";	-- 0x13E0
		when 005089 => D <= "11000001";	-- 0x13E1
		when 005090 => D <= "00001011";	-- 0x13E2
		when 005091 => D <= "01110000";	-- 0x13E3
		when 005092 => D <= "00101011";	-- 0x13E4
		when 005093 => D <= "01110001";	-- 0x13E5
		when 005094 => D <= "11110001";	-- 0x13E6
		when 005095 => D <= "11110101";	-- 0x13E7
		when 005096 => D <= "11001101";	-- 0x13E8
		when 005097 => D <= "11000111";	-- 0x13E9
		when 005098 => D <= "00010100";	-- 0x13EA
		when 005099 => D <= "11110001";	-- 0x13EB
		when 005100 => D <= "00101011";	-- 0x13EC
		when 005101 => D <= "01110111";	-- 0x13ED
		when 005102 => D <= "00101010";	-- 0x13EE
		when 005103 => D <= "00011010";	-- 0x13EF
		when 005104 => D <= "01000000";	-- 0x13F0
		when 005105 => D <= "00100010";	-- 0x13F1
		when 005106 => D <= "00010100";	-- 0x13F2
		when 005107 => D <= "01000000";	-- 0x13F3
		when 005108 => D <= "00101011";	-- 0x13F4
		when 005109 => D <= "00110110";	-- 0x13F5
		when 005110 => D <= "10000000";	-- 0x13F6
		when 005111 => D <= "11001001";	-- 0x13F7
		when 005112 => D <= "00101010";	-- 0x13F8
		when 005113 => D <= "00011100";	-- 0x13F9
		when 005114 => D <= "01000000";	-- 0x13FA
		when 005115 => D <= "00101011";	-- 0x13FB
		when 005116 => D <= "01000110";	-- 0x13FC
		when 005117 => D <= "00101011";	-- 0x13FD
		when 005118 => D <= "01001110";	-- 0x13FE
		when 005119 => D <= "00101011";	-- 0x13FF
		when others => D <= "--------";
		end case;
	end process;
end;
