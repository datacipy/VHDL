library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ROM81hlh is
	port(
		Clk	: in std_logic;
		AIn	: in std_logic_vector(11 downto 0);
		D	: out std_logic_vector(7 downto 0)
	);
end ROM81hlh;

architecture rtl of ROM81hlh is
	signal A	: std_logic_vector(12 downto 0);
begin
	A(9 downto 0) <= AIn(9 downto 0);
	A(12 downto 10) <= "101";
	process (A)
	begin
		case to_integer(unsigned(A)) is
		when 005120 => D <= "01010110";	-- 0x1400
		when 005121 => D <= "00101011";	-- 0x1401
		when 005122 => D <= "01011110";	-- 0x1402
		when 005123 => D <= "00101011";	-- 0x1403
		when 005124 => D <= "01111110";	-- 0x1404
		when 005125 => D <= "00100010";	-- 0x1405
		when 005126 => D <= "00011100";	-- 0x1406
		when 005127 => D <= "01000000";	-- 0x1407
		when 005128 => D <= "11001001";	-- 0x1408
		when 005129 => D <= "11001101";	-- 0x1409
		when 005130 => D <= "00011100";	-- 0x140A
		when 005131 => D <= "00010001";	-- 0x140B
		when 005132 => D <= "11000010";	-- 0x140C
		when 005133 => D <= "10011010";	-- 0x140D
		when 005134 => D <= "00001101";	-- 0x140E
		when 005135 => D <= "11001101";	-- 0x140F
		when 005136 => D <= "10100110";	-- 0x1410
		when 005137 => D <= "00001101";	-- 0x1411
		when 005138 => D <= "00100000";	-- 0x1412
		when 005139 => D <= "00001000";	-- 0x1413
		when 005140 => D <= "11001011";	-- 0x1414
		when 005141 => D <= "10110001";	-- 0x1415
		when 005142 => D <= "11001101";	-- 0x1416
		when 005143 => D <= "10100111";	-- 0x1417
		when 005144 => D <= "00010001";	-- 0x1418
		when 005145 => D <= "11001101";	-- 0x1419
		when 005146 => D <= "00011101";	-- 0x141A
		when 005147 => D <= "00001101";	-- 0x141B
		when 005148 => D <= "00111000";	-- 0x141C
		when 005149 => D <= "00001000";	-- 0x141D
		when 005150 => D <= "11000101";	-- 0x141E
		when 005151 => D <= "11001101";	-- 0x141F
		when 005152 => D <= "11110010";	-- 0x1420
		when 005153 => D <= "00001001";	-- 0x1421
		when 005154 => D <= "11001101";	-- 0x1422
		when 005155 => D <= "01100000";	-- 0x1423
		when 005156 => D <= "00001010";	-- 0x1424
		when 005157 => D <= "11000001";	-- 0x1425
		when 005158 => D <= "11001011";	-- 0x1426
		when 005159 => D <= "11111001";	-- 0x1427
		when 005160 => D <= "00000110";	-- 0x1428
		when 005161 => D <= "00000000";	-- 0x1429
		when 005162 => D <= "11000101";	-- 0x142A
		when 005163 => D <= "00100001";	-- 0x142B
		when 005164 => D <= "00000001";	-- 0x142C
		when 005165 => D <= "00000000";	-- 0x142D
		when 005166 => D <= "11001011";	-- 0x142E
		when 005167 => D <= "01110001";	-- 0x142F
		when 005168 => D <= "00100000";	-- 0x1430
		when 005169 => D <= "00000010";	-- 0x1431
		when 005170 => D <= "00101110";	-- 0x1432
		when 005171 => D <= "00000101";	-- 0x1433
		when 005172 => D <= "11101011";	-- 0x1434
		when 005173 => D <= "11100111";	-- 0x1435
		when 005174 => D <= "00100110";	-- 0x1436
		when 005175 => D <= "01000000";	-- 0x1437
		when 005176 => D <= "11001101";	-- 0x1438
		when 005177 => D <= "11011101";	-- 0x1439
		when 005178 => D <= "00010010";	-- 0x143A
		when 005179 => D <= "11011010";	-- 0x143B
		when 005180 => D <= "00110001";	-- 0x143C
		when 005181 => D <= "00010010";	-- 0x143D
		when 005182 => D <= "11100001";	-- 0x143E
		when 005183 => D <= "11000101";	-- 0x143F
		when 005184 => D <= "00100100";	-- 0x1440
		when 005185 => D <= "11100101";	-- 0x1441
		when 005186 => D <= "01100000";	-- 0x1442
		when 005187 => D <= "01101001";	-- 0x1443
		when 005188 => D <= "11001101";	-- 0x1444
		when 005189 => D <= "00000101";	-- 0x1445
		when 005190 => D <= "00010011";	-- 0x1446
		when 005191 => D <= "11101011";	-- 0x1447
		when 005192 => D <= "11011111";	-- 0x1448
		when 005193 => D <= "11111110";	-- 0x1449
		when 005194 => D <= "00011010";	-- 0x144A
		when 005195 => D <= "00101000";	-- 0x144B
		when 005196 => D <= "11101000";	-- 0x144C
		when 005197 => D <= "11111110";	-- 0x144D
		when 005198 => D <= "00010001";	-- 0x144E
		when 005199 => D <= "00100000";	-- 0x144F
		when 005200 => D <= "10111011";	-- 0x1450
		when 005201 => D <= "11100111";	-- 0x1451
		when 005202 => D <= "11000001";	-- 0x1452
		when 005203 => D <= "01111001";	-- 0x1453
		when 005204 => D <= "01101000";	-- 0x1454
		when 005205 => D <= "00100110";	-- 0x1455
		when 005206 => D <= "00000000";	-- 0x1456
		when 005207 => D <= "00100011";	-- 0x1457
		when 005208 => D <= "00100011";	-- 0x1458
		when 005209 => D <= "00101001";	-- 0x1459
		when 005210 => D <= "00011001";	-- 0x145A
		when 005211 => D <= "11011010";	-- 0x145B
		when 005212 => D <= "11010011";	-- 0x145C
		when 005213 => D <= "00001110";	-- 0x145D
		when 005214 => D <= "11010101";	-- 0x145E
		when 005215 => D <= "11000101";	-- 0x145F
		when 005216 => D <= "11100101";	-- 0x1460
		when 005217 => D <= "01000100";	-- 0x1461
		when 005218 => D <= "01001101";	-- 0x1462
		when 005219 => D <= "00101010";	-- 0x1463
		when 005220 => D <= "00010100";	-- 0x1464
		when 005221 => D <= "01000000";	-- 0x1465
		when 005222 => D <= "00101011";	-- 0x1466
		when 005223 => D <= "11001101";	-- 0x1467
		when 005224 => D <= "10011110";	-- 0x1468
		when 005225 => D <= "00001001";	-- 0x1469
		when 005226 => D <= "00100011";	-- 0x146A
		when 005227 => D <= "01110111";	-- 0x146B
		when 005228 => D <= "11000001";	-- 0x146C
		when 005229 => D <= "00001011";	-- 0x146D
		when 005230 => D <= "00001011";	-- 0x146E
		when 005231 => D <= "00001011";	-- 0x146F
		when 005232 => D <= "00100011";	-- 0x1470
		when 005233 => D <= "01110001";	-- 0x1471
		when 005234 => D <= "00100011";	-- 0x1472
		when 005235 => D <= "01110000";	-- 0x1473
		when 005236 => D <= "11110001";	-- 0x1474
		when 005237 => D <= "00100011";	-- 0x1475
		when 005238 => D <= "01110111";	-- 0x1476
		when 005239 => D <= "01100010";	-- 0x1477
		when 005240 => D <= "01101011";	-- 0x1478
		when 005241 => D <= "00011011";	-- 0x1479
		when 005242 => D <= "00110110";	-- 0x147A
		when 005243 => D <= "00000000";	-- 0x147B
		when 005244 => D <= "11000001";	-- 0x147C
		when 005245 => D <= "11101101";	-- 0x147D
		when 005246 => D <= "10111000";	-- 0x147E
		when 005247 => D <= "11000001";	-- 0x147F
		when 005248 => D <= "01110000";	-- 0x1480
		when 005249 => D <= "00101011";	-- 0x1481
		when 005250 => D <= "01110001";	-- 0x1482
		when 005251 => D <= "00101011";	-- 0x1483
		when 005252 => D <= "00111101";	-- 0x1484
		when 005253 => D <= "00100000";	-- 0x1485
		when 005254 => D <= "11111000";	-- 0x1486
		when 005255 => D <= "11001001";	-- 0x1487
		when 005256 => D <= "00101010";	-- 0x1488
		when 005257 => D <= "00011010";	-- 0x1489
		when 005258 => D <= "01000000";	-- 0x148A
		when 005259 => D <= "00101011";	-- 0x148B
		when 005260 => D <= "11001101";	-- 0x148C
		when 005261 => D <= "10011110";	-- 0x148D
		when 005262 => D <= "00001001";	-- 0x148E
		when 005263 => D <= "00100011";	-- 0x148F
		when 005264 => D <= "00100011";	-- 0x1490
		when 005265 => D <= "11000001";	-- 0x1491
		when 005266 => D <= "11101101";	-- 0x1492
		when 005267 => D <= "01000011";	-- 0x1493
		when 005268 => D <= "00010100";	-- 0x1494
		when 005269 => D <= "01000000";	-- 0x1495
		when 005270 => D <= "11000001";	-- 0x1496
		when 005271 => D <= "11101011";	-- 0x1497
		when 005272 => D <= "00100011";	-- 0x1498
		when 005273 => D <= "11001001";	-- 0x1499
		when 005274 => D <= "00101010";	-- 0x149A
		when 005275 => D <= "00010000";	-- 0x149B
		when 005276 => D <= "01000000";	-- 0x149C
		when 005277 => D <= "00110110";	-- 0x149D
		when 005278 => D <= "10000000";	-- 0x149E
		when 005279 => D <= "00100011";	-- 0x149F
		when 005280 => D <= "00100010";	-- 0x14A0
		when 005281 => D <= "00010100";	-- 0x14A1
		when 005282 => D <= "01000000";	-- 0x14A2
		when 005283 => D <= "00101010";	-- 0x14A3
		when 005284 => D <= "00010100";	-- 0x14A4
		when 005285 => D <= "01000000";	-- 0x14A5
		when 005286 => D <= "00100010";	-- 0x14A6
		when 005287 => D <= "00011010";	-- 0x14A7
		when 005288 => D <= "01000000";	-- 0x14A8
		when 005289 => D <= "00100010";	-- 0x14A9
		when 005290 => D <= "00011100";	-- 0x14AA
		when 005291 => D <= "01000000";	-- 0x14AB
		when 005292 => D <= "11001001";	-- 0x14AC
		when 005293 => D <= "00101010";	-- 0x14AD
		when 005294 => D <= "00010100";	-- 0x14AE
		when 005295 => D <= "01000000";	-- 0x14AF
		when 005296 => D <= "00110110";	-- 0x14B0
		when 005297 => D <= "01111111";	-- 0x14B1
		when 005298 => D <= "00100011";	-- 0x14B2
		when 005299 => D <= "00110110";	-- 0x14B3
		when 005300 => D <= "01110110";	-- 0x14B4
		when 005301 => D <= "00100011";	-- 0x14B5
		when 005302 => D <= "11111101";	-- 0x14B6
		when 005303 => D <= "00110110";	-- 0x14B7
		when 005304 => D <= "00100010";	-- 0x14B8
		when 005305 => D <= "00000010";	-- 0x14B9
		when 005306 => D <= "00011000";	-- 0x14BA
		when 005307 => D <= "11101010";	-- 0x14BB
		when 005308 => D <= "00100001";	-- 0x14BC
		when 005309 => D <= "01011101";	-- 0x14BD
		when 005310 => D <= "01000000";	-- 0x14BE
		when 005311 => D <= "00100010";	-- 0x14BF
		when 005312 => D <= "00011111";	-- 0x14C0
		when 005313 => D <= "01000000";	-- 0x14C1
		when 005314 => D <= "00101010";	-- 0x14C2
		when 005315 => D <= "00011010";	-- 0x14C3
		when 005316 => D <= "01000000";	-- 0x14C4
		when 005317 => D <= "00011000";	-- 0x14C5
		when 005318 => D <= "11100010";	-- 0x14C6
		when 005319 => D <= "11101101";	-- 0x14C7
		when 005320 => D <= "01011011";	-- 0x14C8
		when 005321 => D <= "00010100";	-- 0x14C9
		when 005322 => D <= "01000000";	-- 0x14CA
		when 005323 => D <= "11000011";	-- 0x14CB
		when 005324 => D <= "01011101";	-- 0x14CC
		when 005325 => D <= "00001010";	-- 0x14CD
		when 005326 => D <= "11111110";	-- 0x14CE
		when 005327 => D <= "00100110";	-- 0x14CF
		when 005328 => D <= "00011000";	-- 0x14D0
		when 005329 => D <= "00000010";	-- 0x14D1
		when 005330 => D <= "11111110";	-- 0x14D2
		when 005331 => D <= "00011100";	-- 0x14D3
		when 005332 => D <= "00111111";	-- 0x14D4
		when 005333 => D <= "11010000";	-- 0x14D5
		when 005334 => D <= "11111110";	-- 0x14D6
		when 005335 => D <= "01000000";	-- 0x14D7
		when 005336 => D <= "11001001";	-- 0x14D8
		when 005337 => D <= "11001101";	-- 0x14D9
		when 005338 => D <= "01001000";	-- 0x14DA
		when 005339 => D <= "00010101";	-- 0x14DB
		when 005340 => D <= "11111110";	-- 0x14DC
		when 005341 => D <= "00011011";	-- 0x14DD
		when 005342 => D <= "00100000";	-- 0x14DE
		when 005343 => D <= "00010101";	-- 0x14DF
		when 005344 => D <= "11101111";	-- 0x14E0
		when 005345 => D <= "10100001";	-- 0x14E1
		when 005346 => D <= "11000000";	-- 0x14E2
		when 005347 => D <= "00000010";	-- 0x14E3
		when 005348 => D <= "00110100";	-- 0x14E4
		when 005349 => D <= "11100111";	-- 0x14E5
		when 005350 => D <= "11001101";	-- 0x14E6
		when 005351 => D <= "00010100";	-- 0x14E7
		when 005352 => D <= "00010101";	-- 0x14E8
		when 005353 => D <= "00111000";	-- 0x14E9
		when 005354 => D <= "00001010";	-- 0x14EA
		when 005355 => D <= "11101111";	-- 0x14EB
		when 005356 => D <= "11100000";	-- 0x14EC
		when 005357 => D <= "10100100";	-- 0x14ED
		when 005358 => D <= "00000101";	-- 0x14EE
		when 005359 => D <= "11000000";	-- 0x14EF
		when 005360 => D <= "00000100";	-- 0x14F0
		when 005361 => D <= "00001111";	-- 0x14F1
		when 005362 => D <= "00110100";	-- 0x14F2
		when 005363 => D <= "00011000";	-- 0x14F3
		when 005364 => D <= "11110000";	-- 0x14F4
		when 005365 => D <= "11111110";	-- 0x14F5
		when 005366 => D <= "00101010";	-- 0x14F6
		when 005367 => D <= "11000000";	-- 0x14F7
		when 005368 => D <= "11111101";	-- 0x14F8
		when 005369 => D <= "00110110";	-- 0x14F9
		when 005370 => D <= "01011101";	-- 0x14FA
		when 005371 => D <= "11111111";	-- 0x14FB
		when 005372 => D <= "11100111";	-- 0x14FC
		when 005373 => D <= "11111110";	-- 0x14FD
		when 005374 => D <= "00010101";	-- 0x14FE
		when 005375 => D <= "00101000";	-- 0x14FF
		when 005376 => D <= "00000111";	-- 0x1500
		when 005377 => D <= "11111110";	-- 0x1501
		when 005378 => D <= "00010110";	-- 0x1502
		when 005379 => D <= "00100000";	-- 0x1503
		when 005380 => D <= "00000100";	-- 0x1504
		when 005381 => D <= "11111101";	-- 0x1505
		when 005382 => D <= "00110100";	-- 0x1506
		when 005383 => D <= "01011101";	-- 0x1507
		when 005384 => D <= "11100111";	-- 0x1508
		when 005385 => D <= "11001101";	-- 0x1509
		when 005386 => D <= "01001000";	-- 0x150A
		when 005387 => D <= "00010101";	-- 0x150B
		when 005388 => D <= "11101111";	-- 0x150C
		when 005389 => D <= "11100000";	-- 0x150D
		when 005390 => D <= "00000000";	-- 0x150E
		when 005391 => D <= "00000010";	-- 0x150F
		when 005392 => D <= "00011000";	-- 0x1510
		when 005393 => D <= "00111000";	-- 0x1511
		when 005394 => D <= "00110100";	-- 0x1512
		when 005395 => D <= "11001001";	-- 0x1513
		when 005396 => D <= "11111110";	-- 0x1514
		when 005397 => D <= "00011100";	-- 0x1515
		when 005398 => D <= "11011000";	-- 0x1516
		when 005399 => D <= "11111110";	-- 0x1517
		when 005400 => D <= "00100110";	-- 0x1518
		when 005401 => D <= "00111111";	-- 0x1519
		when 005402 => D <= "11011000";	-- 0x151A
		when 005403 => D <= "11010110";	-- 0x151B
		when 005404 => D <= "00011100";	-- 0x151C
		when 005405 => D <= "01001111";	-- 0x151D
		when 005406 => D <= "00000110";	-- 0x151E
		when 005407 => D <= "00000000";	-- 0x151F
		when 005408 => D <= "11111101";	-- 0x1520
		when 005409 => D <= "00100001";	-- 0x1521
		when 005410 => D <= "00000000";	-- 0x1522
		when 005411 => D <= "01000000";	-- 0x1523
		when 005412 => D <= "11000101";	-- 0x1524
		when 005413 => D <= "11101111";	-- 0x1525
		when 005414 => D <= "10100000";	-- 0x1526
		when 005415 => D <= "00110100";	-- 0x1527
		when 005416 => D <= "11000001";	-- 0x1528
		when 005417 => D <= "00110110";	-- 0x1529
		when 005418 => D <= "10010001";	-- 0x152A
		when 005419 => D <= "01111000";	-- 0x152B
		when 005420 => D <= "10100111";	-- 0x152C
		when 005421 => D <= "00100000";	-- 0x152D
		when 005422 => D <= "00000111";	-- 0x152E
		when 005423 => D <= "01110111";	-- 0x152F
		when 005424 => D <= "10110001";	-- 0x1530
		when 005425 => D <= "11001000";	-- 0x1531
		when 005426 => D <= "01000001";	-- 0x1532
		when 005427 => D <= "01001110";	-- 0x1533
		when 005428 => D <= "00110110";	-- 0x1534
		when 005429 => D <= "10001001";	-- 0x1535
		when 005430 => D <= "00110101";	-- 0x1536
		when 005431 => D <= "11001011";	-- 0x1537
		when 005432 => D <= "00100001";	-- 0x1538
		when 005433 => D <= "11001011";	-- 0x1539
		when 005434 => D <= "00010000";	-- 0x153A
		when 005435 => D <= "00110000";	-- 0x153B
		when 005436 => D <= "11111001";	-- 0x153C
		when 005437 => D <= "11001011";	-- 0x153D
		when 005438 => D <= "00111000";	-- 0x153E
		when 005439 => D <= "11001011";	-- 0x153F
		when 005440 => D <= "00011001";	-- 0x1540
		when 005441 => D <= "00100011";	-- 0x1541
		when 005442 => D <= "01110000";	-- 0x1542
		when 005443 => D <= "00100011";	-- 0x1543
		when 005444 => D <= "01110001";	-- 0x1544
		when 005445 => D <= "00101011";	-- 0x1545
		when 005446 => D <= "00101011";	-- 0x1546
		when 005447 => D <= "11001001";	-- 0x1547
		when 005448 => D <= "11110101";	-- 0x1548
		when 005449 => D <= "11101111";	-- 0x1549
		when 005450 => D <= "10100000";	-- 0x154A
		when 005451 => D <= "00110100";	-- 0x154B
		when 005452 => D <= "11110001";	-- 0x154C
		when 005453 => D <= "11001101";	-- 0x154D
		when 005454 => D <= "00010100";	-- 0x154E
		when 005455 => D <= "00010101";	-- 0x154F
		when 005456 => D <= "11011000";	-- 0x1550
		when 005457 => D <= "11101111";	-- 0x1551
		when 005458 => D <= "00000001";	-- 0x1552
		when 005459 => D <= "10100100";	-- 0x1553
		when 005460 => D <= "00000100";	-- 0x1554
		when 005461 => D <= "00001111";	-- 0x1555
		when 005462 => D <= "00110100";	-- 0x1556
		when 005463 => D <= "11100111";	-- 0x1557
		when 005464 => D <= "00011000";	-- 0x1558
		when 005465 => D <= "11110011";	-- 0x1559
		when 005466 => D <= "11101111";	-- 0x155A
		when 005467 => D <= "00101101";	-- 0x155B
		when 005468 => D <= "00110010";	-- 0x155C
		when 005469 => D <= "11000000";	-- 0x155D
		when 005470 => D <= "00000010";	-- 0x155E
		when 005471 => D <= "00100111";	-- 0x155F
		when 005472 => D <= "10100001";	-- 0x1560
		when 005473 => D <= "00000011";	-- 0x1561
		when 005474 => D <= "00101101";	-- 0x1562
		when 005475 => D <= "00110010";	-- 0x1563
		when 005476 => D <= "00000000";	-- 0x1564
		when 005477 => D <= "00100010";	-- 0x1565
		when 005478 => D <= "00101101";	-- 0x1566
		when 005479 => D <= "00110000";	-- 0x1567
		when 005480 => D <= "00110011";	-- 0x1568
		when 005481 => D <= "01000000";	-- 0x1569
		when 005482 => D <= "00000011";	-- 0x156A
		when 005483 => D <= "00101101";	-- 0x156B
		when 005484 => D <= "00110010";	-- 0x156C
		when 005485 => D <= "00000000";	-- 0x156D
		when 005486 => D <= "00001100";	-- 0x156E
		when 005487 => D <= "00000001";	-- 0x156F
		when 005488 => D <= "00000010";	-- 0x1570
		when 005489 => D <= "00000001";	-- 0x1571
		when 005490 => D <= "00110000";	-- 0x1572
		when 005491 => D <= "10000000";	-- 0x1573
		when 005492 => D <= "01001000";	-- 0x1574
		when 005493 => D <= "00011000";	-- 0x1575
		when 005494 => D <= "10010110";	-- 0x1576
		when 005495 => D <= "10000000";	-- 0x1577
		when 005496 => D <= "00101111";	-- 0x1578
		when 005497 => D <= "00000100";	-- 0x1579
		when 005498 => D <= "00000010";	-- 0x157A
		when 005499 => D <= "00000001";	-- 0x157B
		when 005500 => D <= "10100100";	-- 0x157C
		when 005501 => D <= "11100000";	-- 0x157D
		when 005502 => D <= "00000000";	-- 0x157E
		when 005503 => D <= "00000100";	-- 0x157F
		when 005504 => D <= "00000100";	-- 0x1580
		when 005505 => D <= "00101111";	-- 0x1581
		when 005506 => D <= "00000010";	-- 0x1582
		when 005507 => D <= "00000101";	-- 0x1583
		when 005508 => D <= "00000001";	-- 0x1584
		when 005509 => D <= "00101111";	-- 0x1585
		when 005510 => D <= "11011010";	-- 0x1586
		when 005511 => D <= "00000010";	-- 0x1587
		when 005512 => D <= "00110100";	-- 0x1588
		when 005513 => D <= "11001001";	-- 0x1589
		when 005514 => D <= "11001101";	-- 0x158A
		when 005515 => D <= "11111000";	-- 0x158B
		when 005516 => D <= "00010011";	-- 0x158C
		when 005517 => D <= "10100111";	-- 0x158D
		when 005518 => D <= "00100000";	-- 0x158E
		when 005519 => D <= "00000101";	-- 0x158F
		when 005520 => D <= "01000111";	-- 0x1590
		when 005521 => D <= "01001111";	-- 0x1591
		when 005522 => D <= "11110101";	-- 0x1592
		when 005523 => D <= "00011000";	-- 0x1593
		when 005524 => D <= "00110001";	-- 0x1594
		when 005525 => D <= "01000011";	-- 0x1595
		when 005526 => D <= "01011001";	-- 0x1596
		when 005527 => D <= "01001010";	-- 0x1597
		when 005528 => D <= "11010110";	-- 0x1598
		when 005529 => D <= "10010001";	-- 0x1599
		when 005530 => D <= "00111111";	-- 0x159A
		when 005531 => D <= "11001011";	-- 0x159B
		when 005532 => D <= "01111000";	-- 0x159C
		when 005533 => D <= "11110101";	-- 0x159D
		when 005534 => D <= "11001011";	-- 0x159E
		when 005535 => D <= "11111000";	-- 0x159F
		when 005536 => D <= "00111000";	-- 0x15A0
		when 005537 => D <= "00100100";	-- 0x15A1
		when 005538 => D <= "00111100";	-- 0x15A2
		when 005539 => D <= "11101101";	-- 0x15A3
		when 005540 => D <= "01000100";	-- 0x15A4
		when 005541 => D <= "11111110";	-- 0x15A5
		when 005542 => D <= "00001000";	-- 0x15A6
		when 005543 => D <= "00111000";	-- 0x15A7
		when 005544 => D <= "00000110";	-- 0x15A8
		when 005545 => D <= "01011001";	-- 0x15A9
		when 005546 => D <= "01001000";	-- 0x15AA
		when 005547 => D <= "00000110";	-- 0x15AB
		when 005548 => D <= "00000000";	-- 0x15AC
		when 005549 => D <= "11010110";	-- 0x15AD
		when 005550 => D <= "00001000";	-- 0x15AE
		when 005551 => D <= "10100111";	-- 0x15AF
		when 005552 => D <= "01010111";	-- 0x15B0
		when 005553 => D <= "01111011";	-- 0x15B1
		when 005554 => D <= "00000111";	-- 0x15B2
		when 005555 => D <= "00101000";	-- 0x15B3
		when 005556 => D <= "00000111";	-- 0x15B4
		when 005557 => D <= "11001011";	-- 0x15B5
		when 005558 => D <= "00111000";	-- 0x15B6
		when 005559 => D <= "11001011";	-- 0x15B7
		when 005560 => D <= "00011001";	-- 0x15B8
		when 005561 => D <= "00010101";	-- 0x15B9
		when 005562 => D <= "00100000";	-- 0x15BA
		when 005563 => D <= "11111001";	-- 0x15BB
		when 005564 => D <= "00110000";	-- 0x15BC
		when 005565 => D <= "00001000";	-- 0x15BD
		when 005566 => D <= "00000011";	-- 0x15BE
		when 005567 => D <= "01111000";	-- 0x15BF
		when 005568 => D <= "10110001";	-- 0x15C0
		when 005569 => D <= "00100000";	-- 0x15C1
		when 005570 => D <= "00000011";	-- 0x15C2
		when 005571 => D <= "11110001";	-- 0x15C3
		when 005572 => D <= "00110111";	-- 0x15C4
		when 005573 => D <= "11110101";	-- 0x15C5
		when 005574 => D <= "11000101";	-- 0x15C6
		when 005575 => D <= "11101111";	-- 0x15C7
		when 005576 => D <= "00110100";	-- 0x15C8
		when 005577 => D <= "11000001";	-- 0x15C9
		when 005578 => D <= "11110001";	-- 0x15CA
		when 005579 => D <= "01111001";	-- 0x15CB
		when 005580 => D <= "11001001";	-- 0x15CC
		when 005581 => D <= "11001101";	-- 0x15CD
		when 005582 => D <= "10001010";	-- 0x15CE
		when 005583 => D <= "00010101";	-- 0x15CF
		when 005584 => D <= "11011000";	-- 0x15D0
		when 005585 => D <= "11110101";	-- 0x15D1
		when 005586 => D <= "00000101";	-- 0x15D2
		when 005587 => D <= "00000100";	-- 0x15D3
		when 005588 => D <= "00101000";	-- 0x15D4
		when 005589 => D <= "00000011";	-- 0x15D5
		when 005590 => D <= "11110001";	-- 0x15D6
		when 005591 => D <= "00110111";	-- 0x15D7
		when 005592 => D <= "11001001";	-- 0x15D8
		when 005593 => D <= "11110001";	-- 0x15D9
		when 005594 => D <= "11001001";	-- 0x15DA
		when 005595 => D <= "11101111";	-- 0x15DB
		when 005596 => D <= "00101101";	-- 0x15DC
		when 005597 => D <= "00110010";	-- 0x15DD
		when 005598 => D <= "00000000";	-- 0x15DE
		when 005599 => D <= "00001011";	-- 0x15DF
		when 005600 => D <= "00101101";	-- 0x15E0
		when 005601 => D <= "00110011";	-- 0x15E1
		when 005602 => D <= "00000000";	-- 0x15E2
		when 005603 => D <= "00001101";	-- 0x15E3
		when 005604 => D <= "00000010";	-- 0x15E4
		when 005605 => D <= "00110100";	-- 0x15E5
		when 005606 => D <= "00111110";	-- 0x15E6
		when 005607 => D <= "00011100";	-- 0x15E7
		when 005608 => D <= "11010111";	-- 0x15E8
		when 005609 => D <= "11001001";	-- 0x15E9
		when 005610 => D <= "00100111";	-- 0x15EA
		when 005611 => D <= "00110100";	-- 0x15EB
		when 005612 => D <= "00111110";	-- 0x15EC
		when 005613 => D <= "00010110";	-- 0x15ED
		when 005614 => D <= "11010111";	-- 0x15EE
		when 005615 => D <= "11101111";	-- 0x15EF
		when 005616 => D <= "00110100";	-- 0x15F0
		when 005617 => D <= "01111110";	-- 0x15F1
		when 005618 => D <= "11001101";	-- 0x15F2
		when 005619 => D <= "00011101";	-- 0x15F3
		when 005620 => D <= "00010101";	-- 0x15F4
		when 005621 => D <= "11101111";	-- 0x15F5
		when 005622 => D <= "00110000";	-- 0x15F6
		when 005623 => D <= "01111000";	-- 0x15F7
		when 005624 => D <= "00000000";	-- 0x15F8
		when 005625 => D <= "10000000";	-- 0x15F9
		when 005626 => D <= "00000011";	-- 0x15FA
		when 005627 => D <= "00110000";	-- 0x15FB
		when 005628 => D <= "11101111";	-- 0x15FC
		when 005629 => D <= "00011010";	-- 0x15FD
		when 005630 => D <= "00100000";	-- 0x15FE
		when 005631 => D <= "10011010";	-- 0x15FF
		when 005632 => D <= "10000101";	-- 0x1600
		when 005633 => D <= "00000100";	-- 0x1601
		when 005634 => D <= "00100100";	-- 0x1602
		when 005635 => D <= "11000001";	-- 0x1603
		when 005636 => D <= "00110000";	-- 0x1604
		when 005637 => D <= "00110100";	-- 0x1605
		when 005638 => D <= "00000000";	-- 0x1606
		when 005639 => D <= "00000011";	-- 0x1607
		when 005640 => D <= "00011000";	-- 0x1608
		when 005641 => D <= "00111000";	-- 0x1609
		when 005642 => D <= "10100010";	-- 0x160A
		when 005643 => D <= "00001111";	-- 0x160B
		when 005644 => D <= "00100100";	-- 0x160C
		when 005645 => D <= "00110100";	-- 0x160D
		when 005646 => D <= "00100001";	-- 0x160E
		when 005647 => D <= "01101011";	-- 0x160F
		when 005648 => D <= "01000000";	-- 0x1610
		when 005649 => D <= "00110110";	-- 0x1611
		when 005650 => D <= "10010000";	-- 0x1612
		when 005651 => D <= "00000110";	-- 0x1613
		when 005652 => D <= "00001010";	-- 0x1614
		when 005653 => D <= "00100011";	-- 0x1615
		when 005654 => D <= "11100101";	-- 0x1616
		when 005655 => D <= "11000101";	-- 0x1617
		when 005656 => D <= "11101111";	-- 0x1618
		when 005657 => D <= "10100100";	-- 0x1619
		when 005658 => D <= "00101110";	-- 0x161A
		when 005659 => D <= "00000001";	-- 0x161B
		when 005660 => D <= "00110100";	-- 0x161C
		when 005661 => D <= "11001101";	-- 0x161D
		when 005662 => D <= "11001101";	-- 0x161E
		when 005663 => D <= "00010101";	-- 0x161F
		when 005664 => D <= "11110110";	-- 0x1620
		when 005665 => D <= "10010000";	-- 0x1621
		when 005666 => D <= "11000001";	-- 0x1622
		when 005667 => D <= "11100001";	-- 0x1623
		when 005668 => D <= "01110111";	-- 0x1624
		when 005669 => D <= "00010000";	-- 0x1625
		when 005670 => D <= "11101110";	-- 0x1626
		when 005671 => D <= "00100011";	-- 0x1627
		when 005672 => D <= "00000001";	-- 0x1628
		when 005673 => D <= "00001000";	-- 0x1629
		when 005674 => D <= "00000000";	-- 0x162A
		when 005675 => D <= "11100101";	-- 0x162B
		when 005676 => D <= "00101011";	-- 0x162C
		when 005677 => D <= "01111110";	-- 0x162D
		when 005678 => D <= "11111110";	-- 0x162E
		when 005679 => D <= "10010000";	-- 0x162F
		when 005680 => D <= "00101000";	-- 0x1630
		when 005681 => D <= "11111010";	-- 0x1631
		when 005682 => D <= "11101101";	-- 0x1632
		when 005683 => D <= "01000010";	-- 0x1633
		when 005684 => D <= "11100101";	-- 0x1634
		when 005685 => D <= "01111110";	-- 0x1635
		when 005686 => D <= "11000110";	-- 0x1636
		when 005687 => D <= "01101011";	-- 0x1637
		when 005688 => D <= "11110101";	-- 0x1638
		when 005689 => D <= "11110001";	-- 0x1639
		when 005690 => D <= "00100011";	-- 0x163A
		when 005691 => D <= "01111110";	-- 0x163B
		when 005692 => D <= "11001110";	-- 0x163C
		when 005693 => D <= "00000000";	-- 0x163D
		when 005694 => D <= "00100111";	-- 0x163E
		when 005695 => D <= "11110101";	-- 0x163F
		when 005696 => D <= "11100110";	-- 0x1640
		when 005697 => D <= "00001111";	-- 0x1641
		when 005698 => D <= "01110111";	-- 0x1642
		when 005699 => D <= "11001011";	-- 0x1643
		when 005700 => D <= "11111110";	-- 0x1644
		when 005701 => D <= "00101000";	-- 0x1645
		when 005702 => D <= "11110010";	-- 0x1646
		when 005703 => D <= "11110001";	-- 0x1647
		when 005704 => D <= "11100001";	-- 0x1648
		when 005705 => D <= "00000110";	-- 0x1649
		when 005706 => D <= "00000110";	-- 0x164A
		when 005707 => D <= "00110110";	-- 0x164B
		when 005708 => D <= "10000000";	-- 0x164C
		when 005709 => D <= "00101011";	-- 0x164D
		when 005710 => D <= "00010000";	-- 0x164E
		when 005711 => D <= "11111011";	-- 0x164F
		when 005712 => D <= "11101111";	-- 0x1650
		when 005713 => D <= "00000010";	-- 0x1651
		when 005714 => D <= "11100001";	-- 0x1652
		when 005715 => D <= "00110100";	-- 0x1653
		when 005716 => D <= "11001101";	-- 0x1654
		when 005717 => D <= "11001101";	-- 0x1655
		when 005718 => D <= "00010101";	-- 0x1656
		when 005719 => D <= "00101000";	-- 0x1657
		when 005720 => D <= "00000010";	-- 0x1658
		when 005721 => D <= "11101101";	-- 0x1659
		when 005722 => D <= "01000100";	-- 0x165A
		when 005723 => D <= "01011111";	-- 0x165B
		when 005724 => D <= "00011100";	-- 0x165C
		when 005725 => D <= "00011100";	-- 0x165D
		when 005726 => D <= "11100001";	-- 0x165E
		when 005727 => D <= "00101011";	-- 0x165F
		when 005728 => D <= "00011101";	-- 0x1660
		when 005729 => D <= "01111110";	-- 0x1661
		when 005730 => D <= "11100110";	-- 0x1662
		when 005731 => D <= "00001111";	-- 0x1663
		when 005732 => D <= "00101000";	-- 0x1664
		when 005733 => D <= "11111001";	-- 0x1665
		when 005734 => D <= "01111011";	-- 0x1666
		when 005735 => D <= "11010110";	-- 0x1667
		when 005736 => D <= "00000101";	-- 0x1668
		when 005737 => D <= "11111110";	-- 0x1669
		when 005738 => D <= "00001000";	-- 0x166A
		when 005739 => D <= "11110010";	-- 0x166B
		when 005740 => D <= "10000010";	-- 0x166C
		when 005741 => D <= "00010110";	-- 0x166D
		when 005742 => D <= "11111110";	-- 0x166E
		when 005743 => D <= "11110110";	-- 0x166F
		when 005744 => D <= "11111010";	-- 0x1670
		when 005745 => D <= "10000010";	-- 0x1671
		when 005746 => D <= "00010110";	-- 0x1672
		when 005747 => D <= "11000110";	-- 0x1673
		when 005748 => D <= "00000110";	-- 0x1674
		when 005749 => D <= "00101000";	-- 0x1675
		when 005750 => D <= "01001000";	-- 0x1676
		when 005751 => D <= "11111010";	-- 0x1677
		when 005752 => D <= "10110010";	-- 0x1678
		when 005753 => D <= "00010110";	-- 0x1679
		when 005754 => D <= "01000111";	-- 0x167A
		when 005755 => D <= "11001101";	-- 0x167B
		when 005756 => D <= "11010000";	-- 0x167C
		when 005757 => D <= "00010110";	-- 0x167D
		when 005758 => D <= "00010000";	-- 0x167E
		when 005759 => D <= "11111011";	-- 0x167F
		when 005760 => D <= "00011000";	-- 0x1680
		when 005761 => D <= "01000000";	-- 0x1681
		when 005762 => D <= "01000011";	-- 0x1682
		when 005763 => D <= "11001101";	-- 0x1683
		when 005764 => D <= "11010000";	-- 0x1684
		when 005765 => D <= "00010110";	-- 0x1685
		when 005766 => D <= "11001101";	-- 0x1686
		when 005767 => D <= "11000010";	-- 0x1687
		when 005768 => D <= "00010110";	-- 0x1688
		when 005769 => D <= "00111110";	-- 0x1689
		when 005770 => D <= "00101010";	-- 0x168A
		when 005771 => D <= "11010111";	-- 0x168B
		when 005772 => D <= "01111000";	-- 0x168C
		when 005773 => D <= "10100111";	-- 0x168D
		when 005774 => D <= "11110010";	-- 0x168E
		when 005775 => D <= "10011000";	-- 0x168F
		when 005776 => D <= "00010110";	-- 0x1690
		when 005777 => D <= "11101101";	-- 0x1691
		when 005778 => D <= "01000100";	-- 0x1692
		when 005779 => D <= "01000111";	-- 0x1693
		when 005780 => D <= "00111110";	-- 0x1694
		when 005781 => D <= "00010110";	-- 0x1695
		when 005782 => D <= "00011000";	-- 0x1696
		when 005783 => D <= "00000010";	-- 0x1697
		when 005784 => D <= "00111110";	-- 0x1698
		when 005785 => D <= "00010101";	-- 0x1699
		when 005786 => D <= "11010111";	-- 0x169A
		when 005787 => D <= "01111000";	-- 0x169B
		when 005788 => D <= "00000110";	-- 0x169C
		when 005789 => D <= "11111111";	-- 0x169D
		when 005790 => D <= "00000100";	-- 0x169E
		when 005791 => D <= "11010110";	-- 0x169F
		when 005792 => D <= "00001010";	-- 0x16A0
		when 005793 => D <= "00110000";	-- 0x16A1
		when 005794 => D <= "11111011";	-- 0x16A2
		when 005795 => D <= "11000110";	-- 0x16A3
		when 005796 => D <= "00001010";	-- 0x16A4
		when 005797 => D <= "01001111";	-- 0x16A5
		when 005798 => D <= "01111000";	-- 0x16A6
		when 005799 => D <= "10100111";	-- 0x16A7
		when 005800 => D <= "00101000";	-- 0x16A8
		when 005801 => D <= "00000011";	-- 0x16A9
		when 005802 => D <= "11001101";	-- 0x16AA
		when 005803 => D <= "11101011";	-- 0x16AB
		when 005804 => D <= "00000111";	-- 0x16AC
		when 005805 => D <= "01111001";	-- 0x16AD
		when 005806 => D <= "11001101";	-- 0x16AE
		when 005807 => D <= "11101011";	-- 0x16AF
		when 005808 => D <= "00000111";	-- 0x16B0
		when 005809 => D <= "11001001";	-- 0x16B1
		when 005810 => D <= "11101101";	-- 0x16B2
		when 005811 => D <= "01000100";	-- 0x16B3
		when 005812 => D <= "01000111";	-- 0x16B4
		when 005813 => D <= "00111110";	-- 0x16B5
		when 005814 => D <= "00011011";	-- 0x16B6
		when 005815 => D <= "11010111";	-- 0x16B7
		when 005816 => D <= "00111110";	-- 0x16B8
		when 005817 => D <= "00011100";	-- 0x16B9
		when 005818 => D <= "11010111";	-- 0x16BA
		when 005819 => D <= "00010000";	-- 0x16BB
		when 005820 => D <= "11111101";	-- 0x16BC
		when 005821 => D <= "00011000";	-- 0x16BD
		when 005822 => D <= "00001001";	-- 0x16BE
		when 005823 => D <= "00111110";	-- 0x16BF
		when 005824 => D <= "00011100";	-- 0x16C0
		when 005825 => D <= "11010111";	-- 0x16C1
		when 005826 => D <= "00110101";	-- 0x16C2
		when 005827 => D <= "00110100";	-- 0x16C3
		when 005828 => D <= "11101000";	-- 0x16C4
		when 005829 => D <= "00111110";	-- 0x16C5
		when 005830 => D <= "00011011";	-- 0x16C6
		when 005831 => D <= "11010111";	-- 0x16C7
		when 005832 => D <= "00110101";	-- 0x16C8
		when 005833 => D <= "00110100";	-- 0x16C9
		when 005834 => D <= "11101000";	-- 0x16CA
		when 005835 => D <= "11001101";	-- 0x16CB
		when 005836 => D <= "11010000";	-- 0x16CC
		when 005837 => D <= "00010110";	-- 0x16CD
		when 005838 => D <= "00011000";	-- 0x16CE
		when 005839 => D <= "11111000";	-- 0x16CF
		when 005840 => D <= "01111110";	-- 0x16D0
		when 005841 => D <= "11100110";	-- 0x16D1
		when 005842 => D <= "00001111";	-- 0x16D2
		when 005843 => D <= "11001101";	-- 0x16D3
		when 005844 => D <= "11101011";	-- 0x16D4
		when 005845 => D <= "00000111";	-- 0x16D5
		when 005846 => D <= "00101011";	-- 0x16D6
		when 005847 => D <= "11001001";	-- 0x16D7
		when 005848 => D <= "01111110";	-- 0x16D8
		when 005849 => D <= "00110110";	-- 0x16D9
		when 005850 => D <= "00000000";	-- 0x16DA
		when 005851 => D <= "10100111";	-- 0x16DB
		when 005852 => D <= "11001000";	-- 0x16DC
		when 005853 => D <= "00100011";	-- 0x16DD
		when 005854 => D <= "11001011";	-- 0x16DE
		when 005855 => D <= "01111110";	-- 0x16DF
		when 005856 => D <= "11001011";	-- 0x16E0
		when 005857 => D <= "11111110";	-- 0x16E1
		when 005858 => D <= "00101011";	-- 0x16E2
		when 005859 => D <= "11001000";	-- 0x16E3
		when 005860 => D <= "11000101";	-- 0x16E4
		when 005861 => D <= "00000001";	-- 0x16E5
		when 005862 => D <= "00000101";	-- 0x16E6
		when 005863 => D <= "00000000";	-- 0x16E7
		when 005864 => D <= "00001001";	-- 0x16E8
		when 005865 => D <= "01000001";	-- 0x16E9
		when 005866 => D <= "01001111";	-- 0x16EA
		when 005867 => D <= "00110111";	-- 0x16EB
		when 005868 => D <= "00101011";	-- 0x16EC
		when 005869 => D <= "01111110";	-- 0x16ED
		when 005870 => D <= "00101111";	-- 0x16EE
		when 005871 => D <= "11001110";	-- 0x16EF
		when 005872 => D <= "00000000";	-- 0x16F0
		when 005873 => D <= "01110111";	-- 0x16F1
		when 005874 => D <= "00010000";	-- 0x16F2
		when 005875 => D <= "11111000";	-- 0x16F3
		when 005876 => D <= "01111001";	-- 0x16F4
		when 005877 => D <= "11000001";	-- 0x16F5
		when 005878 => D <= "11001001";	-- 0x16F6
		when 005879 => D <= "11100101";	-- 0x16F7
		when 005880 => D <= "11110101";	-- 0x16F8
		when 005881 => D <= "01001110";	-- 0x16F9
		when 005882 => D <= "00100011";	-- 0x16FA
		when 005883 => D <= "01000110";	-- 0x16FB
		when 005884 => D <= "01110111";	-- 0x16FC
		when 005885 => D <= "00100011";	-- 0x16FD
		when 005886 => D <= "01111001";	-- 0x16FE
		when 005887 => D <= "01001110";	-- 0x16FF
		when 005888 => D <= "11000101";	-- 0x1700
		when 005889 => D <= "00100011";	-- 0x1701
		when 005890 => D <= "01001110";	-- 0x1702
		when 005891 => D <= "00100011";	-- 0x1703
		when 005892 => D <= "01000110";	-- 0x1704
		when 005893 => D <= "11101011";	-- 0x1705
		when 005894 => D <= "01010111";	-- 0x1706
		when 005895 => D <= "01011110";	-- 0x1707
		when 005896 => D <= "11010101";	-- 0x1708
		when 005897 => D <= "00100011";	-- 0x1709
		when 005898 => D <= "01010110";	-- 0x170A
		when 005899 => D <= "00100011";	-- 0x170B
		when 005900 => D <= "01011110";	-- 0x170C
		when 005901 => D <= "11010101";	-- 0x170D
		when 005902 => D <= "11011001";	-- 0x170E
		when 005903 => D <= "11010001";	-- 0x170F
		when 005904 => D <= "11100001";	-- 0x1710
		when 005905 => D <= "11000001";	-- 0x1711
		when 005906 => D <= "11011001";	-- 0x1712
		when 005907 => D <= "00100011";	-- 0x1713
		when 005908 => D <= "01010110";	-- 0x1714
		when 005909 => D <= "00100011";	-- 0x1715
		when 005910 => D <= "01011110";	-- 0x1716
		when 005911 => D <= "11110001";	-- 0x1717
		when 005912 => D <= "11100001";	-- 0x1718
		when 005913 => D <= "11001001";	-- 0x1719
		when 005914 => D <= "10100111";	-- 0x171A
		when 005915 => D <= "11001000";	-- 0x171B
		when 005916 => D <= "11111110";	-- 0x171C
		when 005917 => D <= "00100001";	-- 0x171D
		when 005918 => D <= "00110000";	-- 0x171E
		when 005919 => D <= "00010110";	-- 0x171F
		when 005920 => D <= "11000101";	-- 0x1720
		when 005921 => D <= "01000111";	-- 0x1721
		when 005922 => D <= "11011001";	-- 0x1722
		when 005923 => D <= "11001011";	-- 0x1723
		when 005924 => D <= "00101101";	-- 0x1724
		when 005925 => D <= "11001011";	-- 0x1725
		when 005926 => D <= "00011010";	-- 0x1726
		when 005927 => D <= "11001011";	-- 0x1727
		when 005928 => D <= "00011011";	-- 0x1728
		when 005929 => D <= "11011001";	-- 0x1729
		when 005930 => D <= "11001011";	-- 0x172A
		when 005931 => D <= "00011010";	-- 0x172B
		when 005932 => D <= "11001011";	-- 0x172C
		when 005933 => D <= "00011011";	-- 0x172D
		when 005934 => D <= "00010000";	-- 0x172E
		when 005935 => D <= "11110010";	-- 0x172F
		when 005936 => D <= "11000001";	-- 0x1730
		when 005937 => D <= "11010000";	-- 0x1731
		when 005938 => D <= "11001101";	-- 0x1732
		when 005939 => D <= "01000001";	-- 0x1733
		when 005940 => D <= "00010111";	-- 0x1734
		when 005941 => D <= "11000000";	-- 0x1735
		when 005942 => D <= "11011001";	-- 0x1736
		when 005943 => D <= "10101111";	-- 0x1737
		when 005944 => D <= "00101110";	-- 0x1738
		when 005945 => D <= "00000000";	-- 0x1739
		when 005946 => D <= "01010111";	-- 0x173A
		when 005947 => D <= "01011101";	-- 0x173B
		when 005948 => D <= "11011001";	-- 0x173C
		when 005949 => D <= "00010001";	-- 0x173D
		when 005950 => D <= "00000000";	-- 0x173E
		when 005951 => D <= "00000000";	-- 0x173F
		when 005952 => D <= "11001001";	-- 0x1740
		when 005953 => D <= "00011100";	-- 0x1741
		when 005954 => D <= "11000000";	-- 0x1742
		when 005955 => D <= "00010100";	-- 0x1743
		when 005956 => D <= "11000000";	-- 0x1744
		when 005957 => D <= "11011001";	-- 0x1745
		when 005958 => D <= "00011100";	-- 0x1746
		when 005959 => D <= "00100000";	-- 0x1747
		when 005960 => D <= "00000001";	-- 0x1748
		when 005961 => D <= "00010100";	-- 0x1749
		when 005962 => D <= "11011001";	-- 0x174A
		when 005963 => D <= "11001001";	-- 0x174B
		when 005964 => D <= "00011010";	-- 0x174C
		when 005965 => D <= "10100111";	-- 0x174D
		when 005966 => D <= "11001000";	-- 0x174E
		when 005967 => D <= "00010011";	-- 0x174F
		when 005968 => D <= "00011010";	-- 0x1750
		when 005969 => D <= "11101110";	-- 0x1751
		when 005970 => D <= "10000000";	-- 0x1752
		when 005971 => D <= "00010010";	-- 0x1753
		when 005972 => D <= "00011011";	-- 0x1754
		when 005973 => D <= "11011001";	-- 0x1755
		when 005974 => D <= "11100101";	-- 0x1756
		when 005975 => D <= "11011001";	-- 0x1757
		when 005976 => D <= "11010101";	-- 0x1758
		when 005977 => D <= "11100101";	-- 0x1759
		when 005978 => D <= "11001101";	-- 0x175A
		when 005979 => D <= "11011000";	-- 0x175B
		when 005980 => D <= "00010110";	-- 0x175C
		when 005981 => D <= "01000111";	-- 0x175D
		when 005982 => D <= "11101011";	-- 0x175E
		when 005983 => D <= "11001101";	-- 0x175F
		when 005984 => D <= "11011000";	-- 0x1760
		when 005985 => D <= "00010110";	-- 0x1761
		when 005986 => D <= "01001111";	-- 0x1762
		when 005987 => D <= "10111000";	-- 0x1763
		when 005988 => D <= "00110000";	-- 0x1764
		when 005989 => D <= "00000011";	-- 0x1765
		when 005990 => D <= "01111000";	-- 0x1766
		when 005991 => D <= "01000001";	-- 0x1767
		when 005992 => D <= "11101011";	-- 0x1768
		when 005993 => D <= "11110101";	-- 0x1769
		when 005994 => D <= "10010000";	-- 0x176A
		when 005995 => D <= "11001101";	-- 0x176B
		when 005996 => D <= "11110111";	-- 0x176C
		when 005997 => D <= "00010110";	-- 0x176D
		when 005998 => D <= "11001101";	-- 0x176E
		when 005999 => D <= "00011010";	-- 0x176F
		when 006000 => D <= "00010111";	-- 0x1770
		when 006001 => D <= "11110001";	-- 0x1771
		when 006002 => D <= "11100001";	-- 0x1772
		when 006003 => D <= "01110111";	-- 0x1773
		when 006004 => D <= "11100101";	-- 0x1774
		when 006005 => D <= "01101000";	-- 0x1775
		when 006006 => D <= "01100001";	-- 0x1776
		when 006007 => D <= "00011001";	-- 0x1777
		when 006008 => D <= "11011001";	-- 0x1778
		when 006009 => D <= "11101011";	-- 0x1779
		when 006010 => D <= "11101101";	-- 0x177A
		when 006011 => D <= "01001010";	-- 0x177B
		when 006012 => D <= "11101011";	-- 0x177C
		when 006013 => D <= "01111100";	-- 0x177D
		when 006014 => D <= "10001101";	-- 0x177E
		when 006015 => D <= "01101111";	-- 0x177F
		when 006016 => D <= "00011111";	-- 0x1780
		when 006017 => D <= "10101101";	-- 0x1781
		when 006018 => D <= "11011001";	-- 0x1782
		when 006019 => D <= "11101011";	-- 0x1783
		when 006020 => D <= "11100001";	-- 0x1784
		when 006021 => D <= "00011111";	-- 0x1785
		when 006022 => D <= "00110000";	-- 0x1786
		when 006023 => D <= "00001000";	-- 0x1787
		when 006024 => D <= "00111110";	-- 0x1788
		when 006025 => D <= "00000001";	-- 0x1789
		when 006026 => D <= "11001101";	-- 0x178A
		when 006027 => D <= "00011010";	-- 0x178B
		when 006028 => D <= "00010111";	-- 0x178C
		when 006029 => D <= "00110100";	-- 0x178D
		when 006030 => D <= "00101000";	-- 0x178E
		when 006031 => D <= "00100011";	-- 0x178F
		when 006032 => D <= "11011001";	-- 0x1790
		when 006033 => D <= "01111101";	-- 0x1791
		when 006034 => D <= "11100110";	-- 0x1792
		when 006035 => D <= "10000000";	-- 0x1793
		when 006036 => D <= "11011001";	-- 0x1794
		when 006037 => D <= "00100011";	-- 0x1795
		when 006038 => D <= "01110111";	-- 0x1796
		when 006039 => D <= "00101011";	-- 0x1797
		when 006040 => D <= "00101000";	-- 0x1798
		when 006041 => D <= "00011111";	-- 0x1799
		when 006042 => D <= "01111011";	-- 0x179A
		when 006043 => D <= "11101101";	-- 0x179B
		when 006044 => D <= "01000100";	-- 0x179C
		when 006045 => D <= "00111111";	-- 0x179D
		when 006046 => D <= "01011111";	-- 0x179E
		when 006047 => D <= "01111010";	-- 0x179F
		when 006048 => D <= "00101111";	-- 0x17A0
		when 006049 => D <= "11001110";	-- 0x17A1
		when 006050 => D <= "00000000";	-- 0x17A2
		when 006051 => D <= "01010111";	-- 0x17A3
		when 006052 => D <= "11011001";	-- 0x17A4
		when 006053 => D <= "01111011";	-- 0x17A5
		when 006054 => D <= "00101111";	-- 0x17A6
		when 006055 => D <= "11001110";	-- 0x17A7
		when 006056 => D <= "00000000";	-- 0x17A8
		when 006057 => D <= "01011111";	-- 0x17A9
		when 006058 => D <= "01111010";	-- 0x17AA
		when 006059 => D <= "00101111";	-- 0x17AB
		when 006060 => D <= "11001110";	-- 0x17AC
		when 006061 => D <= "00000000";	-- 0x17AD
		when 006062 => D <= "00110000";	-- 0x17AE
		when 006063 => D <= "00000111";	-- 0x17AF
		when 006064 => D <= "00011111";	-- 0x17B0
		when 006065 => D <= "11011001";	-- 0x17B1
		when 006066 => D <= "00110100";	-- 0x17B2
		when 006067 => D <= "11001010";	-- 0x17B3
		when 006068 => D <= "10000000";	-- 0x17B4
		when 006069 => D <= "00011000";	-- 0x17B5
		when 006070 => D <= "11011001";	-- 0x17B6
		when 006071 => D <= "01010111";	-- 0x17B7
		when 006072 => D <= "11011001";	-- 0x17B8
		when 006073 => D <= "10101111";	-- 0x17B9
		when 006074 => D <= "00011000";	-- 0x17BA
		when 006075 => D <= "01101100";	-- 0x17BB
		when 006076 => D <= "00110111";	-- 0x17BC
		when 006077 => D <= "00110101";	-- 0x17BD
		when 006078 => D <= "00110100";	-- 0x17BE
		when 006079 => D <= "11001000";	-- 0x17BF
		when 006080 => D <= "00100011";	-- 0x17C0
		when 006081 => D <= "10101110";	-- 0x17C1
		when 006082 => D <= "11001011";	-- 0x17C2
		when 006083 => D <= "11111110";	-- 0x17C3
		when 006084 => D <= "00101011";	-- 0x17C4
		when 006085 => D <= "11001001";	-- 0x17C5
		when 006086 => D <= "10101111";	-- 0x17C6
		when 006087 => D <= "11001101";	-- 0x17C7
		when 006088 => D <= "10111100";	-- 0x17C8
		when 006089 => D <= "00010111";	-- 0x17C9
		when 006090 => D <= "11011000";	-- 0x17CA
		when 006091 => D <= "11011001";	-- 0x17CB
		when 006092 => D <= "11100101";	-- 0x17CC
		when 006093 => D <= "11011001";	-- 0x17CD
		when 006094 => D <= "11010101";	-- 0x17CE
		when 006095 => D <= "11101011";	-- 0x17CF
		when 006096 => D <= "11001101";	-- 0x17D0
		when 006097 => D <= "10111100";	-- 0x17D1
		when 006098 => D <= "00010111";	-- 0x17D2
		when 006099 => D <= "11101011";	-- 0x17D3
		when 006100 => D <= "00111000";	-- 0x17D4
		when 006101 => D <= "01011010";	-- 0x17D5
		when 006102 => D <= "11100101";	-- 0x17D6
		when 006103 => D <= "11001101";	-- 0x17D7
		when 006104 => D <= "11110111";	-- 0x17D8
		when 006105 => D <= "00010110";	-- 0x17D9
		when 006106 => D <= "01111000";	-- 0x17DA
		when 006107 => D <= "10100111";	-- 0x17DB
		when 006108 => D <= "11101101";	-- 0x17DC
		when 006109 => D <= "01100010";	-- 0x17DD
		when 006110 => D <= "11011001";	-- 0x17DE
		when 006111 => D <= "11100101";	-- 0x17DF
		when 006112 => D <= "11101101";	-- 0x17E0
		when 006113 => D <= "01100010";	-- 0x17E1
		when 006114 => D <= "11011001";	-- 0x17E2
		when 006115 => D <= "00000110";	-- 0x17E3
		when 006116 => D <= "00100001";	-- 0x17E4
		when 006117 => D <= "00011000";	-- 0x17E5
		when 006118 => D <= "00010001";	-- 0x17E6
		when 006119 => D <= "00110000";	-- 0x17E7
		when 006120 => D <= "00000101";	-- 0x17E8
		when 006121 => D <= "00011001";	-- 0x17E9
		when 006122 => D <= "11011001";	-- 0x17EA
		when 006123 => D <= "11101101";	-- 0x17EB
		when 006124 => D <= "01011010";	-- 0x17EC
		when 006125 => D <= "11011001";	-- 0x17ED
		when 006126 => D <= "11011001";	-- 0x17EE
		when 006127 => D <= "11001011";	-- 0x17EF
		when 006128 => D <= "00011100";	-- 0x17F0
		when 006129 => D <= "11001011";	-- 0x17F1
		when 006130 => D <= "00011101";	-- 0x17F2
		when 006131 => D <= "11011001";	-- 0x17F3
		when 006132 => D <= "11001011";	-- 0x17F4
		when 006133 => D <= "00011100";	-- 0x17F5
		when 006134 => D <= "11001011";	-- 0x17F6
		when 006135 => D <= "00011101";	-- 0x17F7
		when 006136 => D <= "11011001";	-- 0x17F8
		when 006137 => D <= "11001011";	-- 0x17F9
		when 006138 => D <= "00011000";	-- 0x17FA
		when 006139 => D <= "11001011";	-- 0x17FB
		when 006140 => D <= "00011001";	-- 0x17FC
		when 006141 => D <= "11011001";	-- 0x17FD
		when 006142 => D <= "11001011";	-- 0x17FE
		when 006143 => D <= "00011001";	-- 0x17FF
		when others => D <= "--------";
		end case;
	end process;
end;
